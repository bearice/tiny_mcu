//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NZ-LV1QN48C6/I5
//Device: GW1NZ-1
//Created Time: Fri Apr 01 19:01:32 2022

module ARGB_Rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire [27:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h000000003555560900000000000000000000000000000009D02210C000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h000000003543346100000000000000000000000000000090211111D000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000C54333356E00000000000000000000000000000F21000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000E543334456A000000000000000000000000000E210000001B00000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000F544444445490000000000000000000000000B2110000000C00000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000145433444461000000000000000000000000821111100000D00000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000155544345547B00000000000000000000000F21110000000F00000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h000000025554455445530000000000000000000000D211111110000F00000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h00000002555445555456E000000000000000000008221111111000FF00000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000345544456554559000000000000000000003111111111110F00000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000355534334665560000000000000000000C43211222110110E00000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000155445556565556C00000000000000009333222211110110F00000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000E565445556545563A09AB000000000090433221112111110E00000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000B3565443344445570CBEA00000CD0ABE6432211211111110D00000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h000000003455544544444357213CA0009F2EE16643222232222110FB00000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000344544555543456977810ABC15864675422221112211100900000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h00000000354442224466688999A8736679998886433233332211100000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000015544454566779999AAA999AAAAA9987654432322101000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h00000000E55444444688889AAABBBBACCBBBAA9887552211111000E000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0C000000C4664355678989AAABCCDBCDDCCCAA9988755443211100B000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000000B265666767898ABBBBCDDDDDEDCCBBA99876654432211E9000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000C455566767999AACCBCDDEEEEDDDBBAAA987755431111CA000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000D6667778888A99ACCBCEEEEEDDDCCBAAA989877544001E9000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h00000000F66678889999899BCBDEFDEEDDDCCBAAAA988886641010A000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000000146688799999AA9ABADEECEDDDDDCAAAAA9888886521109000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000036778988AA9AA99ABBCEEDDDDCDDCAAAAA998888763111B000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000356888887999A989AABDEDDCCCBCCBAAAAAA98888865221A000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h000000048888989988998889ACEECCDCCBBBBAAAAAA98787876531CA00000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h000002577778877789867778ACEECCCCCBBAAAAAA9999877777753F000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000048987776775568656779BDECBCBCAAAAAA9999888777877651C00000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h00002589875321F0146433568ACDCCCBBAAAA9999877677788877640BA000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h000146789861BCDCBAF2422479BDCCBBA999998740EF247888877653DB000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h000023689873FEDD99AC241369BCDCBBA98886086677926888886553FA000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000267899A844427929D53369BCCCBBA9995B56A866B079988876552D000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h00003689AAA866317E1AA55479ACCBBABAA6B65597559089998876542C000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h000D25789AA87742957BA35569BCCBAABB81995676459399998876542FC00000;
defparam prom_inst_0.INIT_RAM_24 = 256'h000C047899A98754465CA35579BCCBAABB10BB8D8347F7A9998866542E000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0009E15899AAA976766FF26689ACCBAAB923EAAC75808AAAA98775432D900000;
defparam prom_inst_0.INIT_RAM_26 = 256'h000AE036889ABBA88777326689ABCCBAB71461ECC07AAAA9988765442C900000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0007CF2457899AABBB98745799BCBBBAA6348A99AAAAA999988765431D000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h0006AD035578899ABB9976689ACCCCBBA987ABAAAAAAA999877665441C900000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0007ACE26676899AAABA86599ACCCCBBAAAABAAAAAAABAA987666542FA000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h00008ABD046778999ABA85699ABBBBBAAABBBBBAAAAAAA9876776430BA000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h000008ACF34577889AA974578AAAAAAAABBBBBBAA999987667765432C9000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h000007BCF1457778899862467899989AACCBBBAAA998889887654321CA000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000008AC01346677787413577887679BCBBBBBA998877777654232FC0000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h00000079AACF356567761E3677788669BBBBBAAA988776654333330CA0000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h00000008889B03555677BC25666776669BBBAA9987654322222211FC00000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h00000068889AC1455567E8C144454435ABBAA9987654FDCCDF00EFFB90000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h00000008BBCD224675670657F11F995ABBAA9998751FDCBCCDCCCEEC00000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h000007A9877ADE2345673965ADDFC39BBAAA9988863DBBBDEFEEF0DA00000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h00007000008EFCD0F15554F98BB37AAAABA9AA999860EEDCE1210FEB00000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h00000000077BFD1443565664ACC289999888877765520FF11221FFCA00000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000007000898AB1456655672DC47889999988865650FF0F02320D0000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h00000000779A989AC025533552F3457999A98877764FCCDFDEFF0D0000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000877076799AAC0023230D123455877555323211000EEED000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h00000097000688778BFF11222EDF23466766564443E002231BB0000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h000007000008766788ABEDDEEBAC01446566623FE210001110B0000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h00000000007700086798B9BD10CCCCF233310FDFDDF2100EC000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h00000000500006770687AAF33310FCBDCDDCECDBFFE0110DA000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h000000050000758000989A03444420EDACC9ABACD0EE0DE00000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h000000050056600000889BC1343343FEDDBB899CCBDEEDE00000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000005750000067A8A0001343FBAB99899ACBCE00000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h00000000057000000055879CCCBF21EA888989ACDDDF00000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h00000000BFFF113200000000000000000000000000000002C59975A000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h000000009FDDDF1500000000000000000000000000000025997999C000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h00000008FDBBBBF1E00000000000000000000000000000297777775000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000CFDDBBDBF160000000000000000000000000000977777777600000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000EFDDBBBDDFD200000000000000000000000008B777757777A00000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h00000003FDDBBBDDD150000000000000000000000002B9979777777E00000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h00000005FFDBB9BDDD38000000000000000000000004B9977777777000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h00000007DDDBBDDBDFFB0000000000000000000000CB99999977777200000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h00000007DFDBDDDFDDD1E000000000000000000002BBB9999777774200000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h00000009DFDBBDDFFFDFF400000000000000000005DBB9999977777200000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h00000009DFDBBBBBFFFF13000000000000000000AFDBBBBB9977777200000000;
defparam prom_inst_1.INIT_RAM_0B = 256'h00000005DFDBDFFFDFFFF1800000000000000002DFDBBBB99777775200000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000EDFFBBDDDFDDFF1B40246000000000025FDDBB9999997795E00000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h00000008BFFDBBBBBDDDDF3586E4000008A04601FDDB9BB99999995C00000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h00000000BDFDDDBDDDBBDBF175982000207EE511FDBBBBDBBB99994800000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h00000000BBDDBBDDDFDBDF15313514685D3FD131FDBB99999999977400000000;
defparam prom_inst_1.INIT_RAM_10 = 256'h000000009DBDB977BDFFF355577319FF15775331FDBBDDDDB999977000000000;
defparam prom_inst_1.INIT_RAM_11 = 256'h000000005FDBBBDBDFF1155777777777797977531FFDDBBB9979775000000000;
defparam prom_inst_1.INIT_RAM_12 = 256'h00000000EFDBBBDBBF3333577799997BBB99777533FFB9797797770000000000;
defparam prom_inst_1.INIT_RAM_13 = 256'h0A000000CDFFDBDDF133357779BBD9BDDDBB9975553FFDDBB99977A000000000;
defparam prom_inst_1.INIT_RAM_14 = 256'h0000000089FDFDF1F135377999BDDBDDFDBBB97775311FDDB9B9944000000000;
defparam prom_inst_1.INIT_RAM_15 = 256'h00000000ADDDDFFFF155577BB99DDDDFFDBB997775333FFFD9BBB06000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h00000000EFFF111133355559B9BDFDFFDDDBB9777555533FFF99944000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h000000000FFF131155353559B9BDFDDFDDDBB977775555531FB9B74000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h000000005BFF33133555755799BFDBDDDBDDB777775555553FB9B94000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h000000007F1113135735755799BFFDDDBBDDB7777755555531DBB9A000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h00000007DF3333315555535799DFDDDBB9BD977777753355531DD98000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000B11133335333333577BFFBBDBBB999777777533333531FBE400000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h000007DF11111111331111357BDFBBBBB99977777555533333331D4000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000091311FFFF1DDF1FDF115BDDBBBBB9977775555533333533317C00000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h00057B153FD975E15BFB9BDF39BDBBBB9777775553311333555331F784000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h00059D1333F7A8864407B77B159DBB9997757553D724BD35555331FDE6000000;
defparam prom_inst_1.INIT_RAM_20 = 256'h000079D153190A86EE287B59F59BDB9975555178468ACB15555531FD46000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h00005D133551977FAC10CD99F59BBB997775FE264EE049377755331FBE000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h00007D155773DB5D86F24BD9159BB9999771C62E022469577755331F9A000000;
defparam prom_inst_1.INIT_RAM_23 = 256'h000A7B133575DF5FC5D429DDF59BB9779939C442A2248F777755331FB2800000;
defparam prom_inst_1.INIT_RAM_24 = 256'h0006191355773FB559B647DD159BB977999526224006A5977755331FBE000000;
defparam prom_inst_1.INIT_RAM_25 = 256'h0002C5D1557773DBBBBCE7FF357BB99795B92642004D5999975531FDBE400000;
defparam prom_inst_1.INIT_RAM_26 = 256'h0004C19F335799731FF197F15579BB99939F1B866D399997755311FDBC400000;
defparam prom_inst_1.INIT_RAM_27 = 256'h000E807BD135577997531BD1579B999971DF377799999777755311FD9C000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h000C4A37DF13357797551FF377BBBB997553999999999777553111FD9C400000;
defparam prom_inst_1.INIT_RAM_29 = 256'h000E48C7DF11355797973FF579BBBB99979999999979B977531131D926000000;
defparam prom_inst_1.INIT_RAM_2A = 256'h0000048C39D1135577973DF57999B997979999999779777533331FB7A4000000;
defparam prom_inst_1.INIT_RAM_2B = 256'h0000004A07BD135557751BF35799979779B99999977775313331FDB9C4000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h0000006805BD11133553F9D1357755579BB9BB9977755575331FDDB7C4000000;
defparam prom_inst_1.INIT_RAM_2D = 256'h00000004A139BFF11131B5BF133533359B9999B97755333331FDBB92A0000000;
defparam prom_inst_1.INIT_RAM_2E = 256'h000000E446807DFDF11F509F11133115BB9999997553311FDBBBBB7C60000000;
defparam prom_inst_1.INIT_RAM_2F = 256'h00000000222637DDDF11AC7DFFF111F159997777531FDB997999972C00000000;
defparam prom_inst_1.INIT_RAM_30 = 256'h000000E22244A5BDDDF3E2C7BBDDDBBF9999775531FB2ECCE255222A40000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000068AC77BFFDF13EA025528CF7B97755553F70EAACCECCC02A00000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h000000420004AE79BDF1B6EC8EE00D79977775353FBEA8AC002025E600000000;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000E000002C0AC303BDDB2448A91797797577755315EECC0797720800000000;
defparam prom_inst_1.INIT_RAM_34 = 256'h000000000006EC39B9DFDFFB8AA9355553333131FFF93027799722C600000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h00000000000224639DFFDDF19CCB135557753331FFD5225239B95E0000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h00000000EE244224815DD99DD709BF15777753113FB2ACE202225E0000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h00000000000EE0424681379791C579BDF311FDDB99755353002E000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000002E000C00E006EE35777EC279BF111FFFDDB9E5579B7AA0000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000EE02048CACCC64835BBFDFFF7B2E755557755A0000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000E020628E53AAAA07999530C2CE077730A000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h00000000A0000E000E20440999530C8C8CCAE8C80003773E8000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000C00000C2000202619BBBB75EC6A82486AC3E03E000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000C00CEE000000028859BB9B90EAA86244AC8EE0E000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000CEC00000EE42613339B90848442446C8CE00000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h000000000CE0000000AC0E28A88055E62224246AEEE200000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h00000000A666B7A90000000000000000000000000000000D12AEA2D000000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h00000000A66226B2000000000000000000000000000000D2EAAAAA5000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000000966222E6B100000000000000000000000000000EEAAAAAA6000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h00000001622EEEE6750000000000000000000000000006EAAAAAAAA900000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h00000005662EEE226ED00000000000000000000000009EEAAAAAAAAD00000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000000E662EEE2E2BE000000000000000000000000DEEEAAAAAAAA900000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h000000026622EEE222B5000000000000000000000002EEEAAAAAAAAE00000000;
defparam prom_inst_2.INIT_RAM_07 = 256'h000000066622E22E266A000000000000000000000012EEEEEAAAAAA200000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h00000006662EEE22226B100000000000000000000DE22EEEAAAAAAA200000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h0000000A6622EE2226262D00000000000000000002622EEEEEEEEEA200000000;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000A662EEEEE6666BE000000000000000000D6622222EEEEEEA200000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h00000002662E222626666B90000000000000000D2662222EEEEEEEA200000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h00000005666EEE2262266BA10DD10000000000D2A6622EEE2EEEEEAD00000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h000000092662EEEEE22266BE911D000005D0D5ABA662222EEEEEEEA500000000;
defparam prom_inst_2.INIT_RAM_0E = 256'h0000000022622EE2E22222AB2E69D000D62112BFA662226222EEEEAD00000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h00000000E2662E22222E26BFB7BE6D15EEB2EBFFA6622E2E2EEE2EE500000000;
defparam prom_inst_2.INIT_RAM_10 = 256'h00000000A6262EAAE2666BFFF33B76667F33FFFFA662666222222EE000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h000000002662222E2667BFF333733333373733FFBA66622222222EA000000000;
defparam prom_inst_2.INIT_RAM_12 = 256'h000000005662222EE6BBBB333777777BBB77773FFB6622E2E2222E2000000000;
defparam prom_inst_2.INIT_RAM_13 = 256'h0D000000D2662E2267BFBF3737BBFBBBFBBB7733FFF6A66222222ED000000000;
defparam prom_inst_2.INIT_RAM_14 = 256'h00000000DE62662727BFF377B7BFFBBFFFBBB73333FBB66662222A5000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h00000000D222266627FFF33BB77FFFFFFFBB773373FFF6A66222265000000000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0000000056627777BBBFFF37B7BFFFFFFFFBBB377333FFFAA6222A1000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h00000000A2667B7BFFFFFFF7B7BFFFFFBFFBB7777333FFFBB6622E5000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h000000002E22BB7BFFFF3FF377BFFBFFBBFFB7773333FFFFBA626E5000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0000000062777BBBF3FF3FF377BFFFFFFBFFB7737733FFFFFB666E1000000000;
defparam prom_inst_2.INIT_RAM_1A = 256'h00000006E2BBBBB7FFFFFBF377FFFFFBBBBFB7737773FFFFFBB66E9000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000A777BFBFFBBBFBBF33BFFFBFBBBBBB7737733FFFFFFBB625100000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h000002E2777B7777BBB777BF3BFFFBBBBB77777773333FFFFFFFB22000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h00000A7BB766267226B2E2BB3BFFFBBBBB777773333FFFFFFFFFB7A100000000;
defparam prom_inst_2.INIT_RAM_1E = 256'h000E2A7FB62EA69E2E2EAE26F7BFFFBBB77777373FFFFFF33FFFFB6691000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h00026E7BBB6A11955926E6AEB3BFBBBBB777733FA2EE6E3333FFFB6E55000000;
defparam prom_inst_2.INIT_RAM_20 = 256'h000026E7FF722D5104116E2A63BFFBBB73333F65DDD15E77333FFB6225000000;
defparam prom_inst_2.INIT_RAM_21 = 256'h00002E7BBF3B6EE948295EA66FBBBBB77773A99DD59E2A777733FBB6E5000000;
defparam prom_inst_2.INIT_RAM_22 = 256'h00002E7F337FE6A509595EEA7F7FBB77777F5DE19AE2AA777733FFB6ED000000;
defparam prom_inst_2.INIT_RAM_23 = 256'h00092E7BF3732AA9822D1A2E63BBFB77BB3692268A22AEBB7733FFB6EE900000;
defparam prom_inst_2.INIT_RAM_24 = 256'h0005667BFF33FE2A2AE15A22BFBBBB77BB6EE6AE1EE6A7BB7333FBB6E5000000;
defparam prom_inst_2.INIT_RAM_25 = 256'h00091EEBF3337FE62221DA22B37BFB7773A6E626A26E7BBBB73FFB62E5100000;
defparam prom_inst_2.INIT_RAM_26 = 256'h0001DA62BBF3777F322BEA27F37BFBB7B3AE3A666E7BBBB7333FB762A1100000;
defparam prom_inst_2.INIT_RAM_27 = 256'h00049A6E27BF337777FBBE2B37BFBBB77FE23B77BBBBB77333FBBB62A1000000;
defparam prom_inst_2.INIT_RAM_28 = 256'h00001DE6E27BFF37773FB26F77FFFFB77773BBBBBBBB77733FBBBB62A1100000;
defparam prom_inst_2.INIT_RAM_29 = 256'h00001912E277BF377373B2637BFFFFB777BBBBBBBB7BBB733FBBB72AE5000000;
defparam prom_inst_2.INIT_RAM_2A = 256'h00005151EA277FFF3373B2A37BFFFBB777BBBBBBB77B7733FBBBB2E2D1000000;
defparam prom_inst_2.INIT_RAM_2B = 256'h0000091DA6E27BFFF33F72A37BBFBBB77BBBBBBB777333FBBFFB62EA11000000;
defparam prom_inst_2.INIT_RAM_2C = 256'h000005196EA27B7FBFFB2EA37BBBB7777BFBBBBB7733FF33FB722EE615000000;
defparam prom_inst_2.INIT_RAM_2D = 256'h0000009D9AE6A26777B7EEA277BBB777BBBBBBBB733FFBBBB72EEEAED0000000;
defparam prom_inst_2.INIT_RAM_2E = 256'h0000004D119A6E2227726A6E77777737BBBBB7773FFBB7722EEEEE6150000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h00000009D9D5E6EEE277D56E266773237BB77773FFB62EAA6AAA66E100000000;
defparam prom_inst_2.INIT_RAM_30 = 256'h000000099DD19EAEEE271D1AE22222EEBB773333FB6EE5155EE2AEED10000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h00000009559D22A22E2724C5AAAA552BBB773F33F26A5DD115111AED00000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h000005D95991D126AE23A58CD1566EBBB77333FFF6A5D9D16AAAE25500000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h00000000009169DAAEAEEE6D5916F7B77733333FFF7E5511A2662EA900000000;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000005511DA6A6E2E22219D6F333FFFBFBBB6226EAA26AA6EE1500000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h00000050009D9D5A6A22EE27E596BFF33333FFB726EEEA2EEAEA250000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h00000000449DD9D15A2EEAAE2A6EE6BF3333FF7BB2EAD15EAEEE250000000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h00000009550445DD119AA266A296AEE22BB7222E66622E2EAAA5000000000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h00000090000059459515E226699E6AE2777222EEE65E266A2DD0000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h000005000005500599155D155D91E2EE622226AA52222E2222D0000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h000000000055000949D951952E5511A6AAA2EA1A15A622EA1000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h000000008000005504D9D1A6AA62E5D1911D1915A6AE22E59000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000C00001C9000D9D1A6EEEE62515D9D1959DE5AE5600000000000000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000C00C000000099D99E6EAAEAA5DD9591191955A5A00000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000C0C00000041D1AAAEAA6A91511D115191500000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h000000000C000000008C94D9D99A2E55D991D151555E00000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[27:0],dout[15:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 4;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h00000000DEEEEECA0000000000000000000000000000000ACDDDDDB000000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h00000000DEEEEEED000000000000000000000000000000ADDDDDDDC000000000;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000000BEEEEEDEEC00000000000000000000000000000CDDDDDDDD000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0000000CEEEDDDDEEB000000000000000000000000000CDDDDDDDDDB00000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h0000000CEEEDDDEEEDA0000000000000000000000000BDDDDDDDDDDB00000000;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000000CEEEDDDEDEEC000000000000000000000000ADDDDDDDDDDDC00000000;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000DEEEEDDDEEEEB00000000000000000000000DDDDDDDDDDDDC00000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000000DEEEEDEEDEEED0000000000000000000000CEDDDDDDDDDDDD00000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000DEEEDDDEEEEEEC00000000000000000000ADEEDDDDDDDDDDD00000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000000DEEEEDDEEEEEEEA0000000000000000000DEEEDDDDDDDDDDD00000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000000DEEEDDDDDEEEEEC000000000000000000BEEEEEEEDDDDDDDD00000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000000DEEEDEEEEEEEEEEB0000000000000000AEEEEEEEDDDDDDDDD00000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000000CEEEDDDEEEEEEEEDB0AAB0000000000ADEEEEEDDDEDDDDDDC00000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000000BEEEEDDDDDEEEEEECBBCA00000BB0ABCEEEEEEEEDDDDDDDDC00000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h00000000EEEEEDDEDEEEEEEEDCDBA000ACDCCDEEEEEEEEEEEEDDDDDB00000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h00000000DEEEEDEEEEEDEEEEEEECCABBCDEEDEEEEEEEEDEDEDDDEDDB00000000;
defparam prom_inst_3.INIT_RAM_10 = 256'h00000000DEEEEDDDDEEEEEEEEFFEEDEEEEFFEEEEEEEEEEEEEEEEEDD000000000;
defparam prom_inst_3.INIT_RAM_11 = 256'h00000000DEEEEEEDEEEEEEEFFFFFFFFFFFFFFFEEEEEEEEEEEEEEEDD000000000;
defparam prom_inst_3.INIT_RAM_12 = 256'h00000000CEEEEEEDDEEEEEFFFFFFFFFFFFFFFFFEEEEEEEDEDEEEEDD000000000;
defparam prom_inst_3.INIT_RAM_13 = 256'h0B000000BEEEEDEEEEEEEEFFFFFFFFFFFFFFFFFFEEEEEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h00000000BDEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h00000000BEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h00000000CEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h00000000CEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h00000000DDEEEEEEEEEEFEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h00000000DEEEEEEEEFEEFEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEDC000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000000DDEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEDB000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h0000000DEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEEECB00000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h00000DDEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFFFFFFFFFEEEEEEEEED000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h00000DEEEEEEEEEEEEEEDEEEFFFFFFFFFFFFFFFFFFFEEEEEEEEEEEDC00000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h000CDDEEEEEDDDCCDDEDDDEEEFFFFFFFFFFFFFFFFEEEEEEFFEEEEEEDBB000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h000DDDEEEEEDDCBBBBDDDDDDEFFFFFFFFFFFFFFEEEDDEEFFFFEEEEEDCB000000;
defparam prom_inst_3.INIT_RAM_20 = 256'h0000DDDEEEEEDBBBAABCDDDDEFFFFFFFFFFFFEEDCCCDDEFFFFFEEEEEDB000000;
defparam prom_inst_3.INIT_RAM_21 = 256'h0000DDEEEEFEDCCB99CACDDDEEFFFFFFFFFFEDCCADDDEEFFFFFFEEEEDC000000;
defparam prom_inst_3.INIT_RAM_22 = 256'h0000DDEEFFFEDDCB9ABABDDDEEFFFFFFFFFEDCDDADDEEEFFFFFFEEEEDB000000;
defparam prom_inst_3.INIT_RAM_23 = 256'h000BDDEEEFFFEDCB9CDABDEDEFFFFFFFFFFEDEED9DEEEEFFFFFFEEEEDCB00000;
defparam prom_inst_3.INIT_RAM_24 = 256'h000BCDEEEEFFEDDCCCCBBDEEEEFFFFFFFFEDDEDCBDDEEFFFFFFFEEEEDC000000;
defparam prom_inst_3.INIT_RAM_25 = 256'h000ACCDEEFFFFEDDDDDCCDEEEFFFFFFFFFEEDEEDDEEEFFFFFFFEEEEEDCB00000;
defparam prom_inst_3.INIT_RAM_26 = 256'h000BBCDEEEEFFFFEEEEEDDEEEFFFFFFFFFEEFEEEEEFFFFFFFFFEEEEEDCB00000;
defparam prom_inst_3.INIT_RAM_27 = 256'h000ABCDDEEEEFFFFFFEEEDEEFFFFFFFFFEEFFFFFFFFFFFFFFFEEEEEEDC000000;
defparam prom_inst_3.INIT_RAM_28 = 256'h000ABBCDDEEEEEFFFFFEEEEEFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEDCB00000;
defparam prom_inst_3.INIT_RAM_29 = 256'h000ABBCDDEEEEEFFFFFFEEEFFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEDCB000000;
defparam prom_inst_3.INIT_RAM_2A = 256'h0000ABBCCDEEEEEEFFFFEEEFFFFFFFFFFFFFFFFFFFFFFFFFEEEEEEDDBB000000;
defparam prom_inst_3.INIT_RAM_2B = 256'h00000ABBCDDEEEEEEFFEEEEFFFFFFFFFFFFFFFFFFFFFFFEEEEEEEEDDCB000000;
defparam prom_inst_3.INIT_RAM_2C = 256'h00000ABBCCDEEEEEEEEEEDEFFFFFFFFFFFFFFFFFFFFFEEFFEEEEEDDDCB000000;
defparam prom_inst_3.INIT_RAM_2D = 256'h000000AABCCDDEEEEEEEDDEFFFFFFFFFFFFFFFFFFFFEEEEEEEEDDDDCB0000000;
defparam prom_inst_3.INIT_RAM_2E = 256'h000000AABBBCDDEEEEEEDDEEFFFFFFFFFFFFFFFFFEEEEEEEEDDDDDDCB0000000;
defparam prom_inst_3.INIT_RAM_2F = 256'h0000000AAAABCDDDDEEECDEEFFFFFFFFFFFFFFFFEEEEEDDDDDDDDDCC00000000;
defparam prom_inst_3.INIT_RAM_30 = 256'h000000AAAAABBCDDDDEEDCEEEFFFFFEEFFFFFFFFEEEDCCCCCCCDCCCBB0000000;
defparam prom_inst_3.INIT_RAM_31 = 256'h0000000ABBBBDDDEEDEEDCCDEEEEEEFFFFFFFEFFEEDCCBBCCCCCCCCB00000000;
defparam prom_inst_3.INIT_RAM_32 = 256'h00000AAAAAABBCDDDDEEDCCCDEEEEEFFFFFFFFEEEEDCBBBCCCCCCDCB00000000;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000A00000ACCBBCCCDDDDDCDDEEEFFFFFFFFFFEEEECCCCCCDDDDCCB00000000;
defparam prom_inst_3.INIT_RAM_34 = 256'h000000000AABCBCDDDDEDEEEDDDEEFFFEEEEEEEEEEEDCCCDDDDDCCCB00000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h000000A000AAAABCDDEEDDEEDDDEEEEFFFFFEEEEEEDCCCDCCDDDDC0000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h00000000AAAAAAABBCDDDDDDEDDDDEEEFFFFEEEEEEDCBCCCCCCCDC0000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000AAA0AAAAABBBCCDDDDDCDDDDEEEEEEEEDDDDDDCDCCCCC000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h000000AA000AAAAAABCCCDDDDCCCDDDEEEEEEEDDDDCCDDDDDBB0000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h00000A00000AAAAAAABBCBCCCBBCCDDDEEEEEDDCCDDDDCDDDDB0000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000AA000AAAAABBBCDCCCCCCDDDDDCCCCCCCDDDCCC000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000090000AAA0AAAABCDDDDDCCBCBCCBCBCBCCCCDDCCB000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h000000090000A9A000AAABCDDDDDDDCCBBBABBBBBCCCCCC00000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h00000009009AA00000AAABBCDDDDDDCCBBBBABBBCBCCCCC00000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h00000000009A900000AABABCCCCDDDCBBBBBABBBCBCC00000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000009A000000099AAABBBBCDCCBAAABABBCCCCC00000000000000000000;

endmodule //ARGB_Rom
