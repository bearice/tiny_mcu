//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NZ-LV1QN48C6/I5
//Device: GW1NZ-1
//Created Time: Fri Apr 01 14:18:16 2022

module Gowin_ROM16 (dout, ad);

output [15:0] dout;
input [7:0] ad;

wire [0:0] rom16_inst_0_dout;
wire [1:1] rom16_inst_1_dout;
wire [2:2] rom16_inst_2_dout;
wire [3:3] rom16_inst_3_dout;
wire [4:4] rom16_inst_4_dout;
wire [5:5] rom16_inst_5_dout;
wire [6:6] rom16_inst_6_dout;
wire [7:7] rom16_inst_7_dout;
wire [8:8] rom16_inst_8_dout;
wire [9:9] rom16_inst_9_dout;
wire [10:10] rom16_inst_10_dout;
wire [11:11] rom16_inst_11_dout;
wire [12:12] rom16_inst_12_dout;
wire [13:13] rom16_inst_13_dout;
wire [14:14] rom16_inst_14_dout;
wire [15:15] rom16_inst_15_dout;
wire [0:0] rom16_inst_16_dout;
wire [1:1] rom16_inst_17_dout;
wire [2:2] rom16_inst_18_dout;
wire [3:3] rom16_inst_19_dout;
wire [4:4] rom16_inst_20_dout;
wire [5:5] rom16_inst_21_dout;
wire [6:6] rom16_inst_22_dout;
wire [7:7] rom16_inst_23_dout;
wire [8:8] rom16_inst_24_dout;
wire [9:9] rom16_inst_25_dout;
wire [10:10] rom16_inst_26_dout;
wire [11:11] rom16_inst_27_dout;
wire [12:12] rom16_inst_28_dout;
wire [13:13] rom16_inst_29_dout;
wire [14:14] rom16_inst_30_dout;
wire [15:15] rom16_inst_31_dout;
wire [0:0] rom16_inst_32_dout;
wire [1:1] rom16_inst_33_dout;
wire [2:2] rom16_inst_34_dout;
wire [3:3] rom16_inst_35_dout;
wire [4:4] rom16_inst_36_dout;
wire [5:5] rom16_inst_37_dout;
wire [6:6] rom16_inst_38_dout;
wire [7:7] rom16_inst_39_dout;
wire [8:8] rom16_inst_40_dout;
wire [9:9] rom16_inst_41_dout;
wire [10:10] rom16_inst_42_dout;
wire [11:11] rom16_inst_43_dout;
wire [12:12] rom16_inst_44_dout;
wire [13:13] rom16_inst_45_dout;
wire [14:14] rom16_inst_46_dout;
wire [15:15] rom16_inst_47_dout;
wire [0:0] rom16_inst_48_dout;
wire [1:1] rom16_inst_49_dout;
wire [2:2] rom16_inst_50_dout;
wire [3:3] rom16_inst_51_dout;
wire [4:4] rom16_inst_52_dout;
wire [5:5] rom16_inst_53_dout;
wire [6:6] rom16_inst_54_dout;
wire [7:7] rom16_inst_55_dout;
wire [8:8] rom16_inst_56_dout;
wire [9:9] rom16_inst_57_dout;
wire [10:10] rom16_inst_58_dout;
wire [11:11] rom16_inst_59_dout;
wire [12:12] rom16_inst_60_dout;
wire [13:13] rom16_inst_61_dout;
wire [14:14] rom16_inst_62_dout;
wire [15:15] rom16_inst_63_dout;
wire [0:0] rom16_inst_64_dout;
wire [1:1] rom16_inst_65_dout;
wire [2:2] rom16_inst_66_dout;
wire [3:3] rom16_inst_67_dout;
wire [4:4] rom16_inst_68_dout;
wire [5:5] rom16_inst_69_dout;
wire [6:6] rom16_inst_70_dout;
wire [7:7] rom16_inst_71_dout;
wire [8:8] rom16_inst_72_dout;
wire [9:9] rom16_inst_73_dout;
wire [10:10] rom16_inst_74_dout;
wire [11:11] rom16_inst_75_dout;
wire [12:12] rom16_inst_76_dout;
wire [13:13] rom16_inst_77_dout;
wire [14:14] rom16_inst_78_dout;
wire [15:15] rom16_inst_79_dout;
wire [0:0] rom16_inst_80_dout;
wire [1:1] rom16_inst_81_dout;
wire [2:2] rom16_inst_82_dout;
wire [3:3] rom16_inst_83_dout;
wire [4:4] rom16_inst_84_dout;
wire [5:5] rom16_inst_85_dout;
wire [6:6] rom16_inst_86_dout;
wire [7:7] rom16_inst_87_dout;
wire [8:8] rom16_inst_88_dout;
wire [9:9] rom16_inst_89_dout;
wire [10:10] rom16_inst_90_dout;
wire [11:11] rom16_inst_91_dout;
wire [12:12] rom16_inst_92_dout;
wire [13:13] rom16_inst_93_dout;
wire [14:14] rom16_inst_94_dout;
wire [15:15] rom16_inst_95_dout;
wire [0:0] rom16_inst_96_dout;
wire [1:1] rom16_inst_97_dout;
wire [2:2] rom16_inst_98_dout;
wire [3:3] rom16_inst_99_dout;
wire [4:4] rom16_inst_100_dout;
wire [5:5] rom16_inst_101_dout;
wire [6:6] rom16_inst_102_dout;
wire [7:7] rom16_inst_103_dout;
wire [8:8] rom16_inst_104_dout;
wire [9:9] rom16_inst_105_dout;
wire [10:10] rom16_inst_106_dout;
wire [11:11] rom16_inst_107_dout;
wire [12:12] rom16_inst_108_dout;
wire [13:13] rom16_inst_109_dout;
wire [14:14] rom16_inst_110_dout;
wire [15:15] rom16_inst_111_dout;
wire [0:0] rom16_inst_112_dout;
wire [1:1] rom16_inst_113_dout;
wire [2:2] rom16_inst_114_dout;
wire [3:3] rom16_inst_115_dout;
wire [4:4] rom16_inst_116_dout;
wire [5:5] rom16_inst_117_dout;
wire [6:6] rom16_inst_118_dout;
wire [7:7] rom16_inst_119_dout;
wire [8:8] rom16_inst_120_dout;
wire [9:9] rom16_inst_121_dout;
wire [10:10] rom16_inst_122_dout;
wire [11:11] rom16_inst_123_dout;
wire [12:12] rom16_inst_124_dout;
wire [13:13] rom16_inst_125_dout;
wire [14:14] rom16_inst_126_dout;
wire [15:15] rom16_inst_127_dout;
wire [0:0] rom16_inst_128_dout;
wire [1:1] rom16_inst_129_dout;
wire [2:2] rom16_inst_130_dout;
wire [3:3] rom16_inst_131_dout;
wire [4:4] rom16_inst_132_dout;
wire [5:5] rom16_inst_133_dout;
wire [6:6] rom16_inst_134_dout;
wire [7:7] rom16_inst_135_dout;
wire [8:8] rom16_inst_136_dout;
wire [9:9] rom16_inst_137_dout;
wire [10:10] rom16_inst_138_dout;
wire [11:11] rom16_inst_139_dout;
wire [12:12] rom16_inst_140_dout;
wire [13:13] rom16_inst_141_dout;
wire [14:14] rom16_inst_142_dout;
wire [15:15] rom16_inst_143_dout;
wire [0:0] rom16_inst_144_dout;
wire [1:1] rom16_inst_145_dout;
wire [2:2] rom16_inst_146_dout;
wire [3:3] rom16_inst_147_dout;
wire [4:4] rom16_inst_148_dout;
wire [5:5] rom16_inst_149_dout;
wire [6:6] rom16_inst_150_dout;
wire [7:7] rom16_inst_151_dout;
wire [8:8] rom16_inst_152_dout;
wire [9:9] rom16_inst_153_dout;
wire [10:10] rom16_inst_154_dout;
wire [11:11] rom16_inst_155_dout;
wire [12:12] rom16_inst_156_dout;
wire [13:13] rom16_inst_157_dout;
wire [14:14] rom16_inst_158_dout;
wire [15:15] rom16_inst_159_dout;
wire [0:0] rom16_inst_160_dout;
wire [1:1] rom16_inst_161_dout;
wire [2:2] rom16_inst_162_dout;
wire [3:3] rom16_inst_163_dout;
wire [4:4] rom16_inst_164_dout;
wire [5:5] rom16_inst_165_dout;
wire [6:6] rom16_inst_166_dout;
wire [7:7] rom16_inst_167_dout;
wire [8:8] rom16_inst_168_dout;
wire [9:9] rom16_inst_169_dout;
wire [10:10] rom16_inst_170_dout;
wire [11:11] rom16_inst_171_dout;
wire [12:12] rom16_inst_172_dout;
wire [13:13] rom16_inst_173_dout;
wire [14:14] rom16_inst_174_dout;
wire [15:15] rom16_inst_175_dout;
wire [0:0] rom16_inst_176_dout;
wire [1:1] rom16_inst_177_dout;
wire [2:2] rom16_inst_178_dout;
wire [3:3] rom16_inst_179_dout;
wire [4:4] rom16_inst_180_dout;
wire [5:5] rom16_inst_181_dout;
wire [6:6] rom16_inst_182_dout;
wire [7:7] rom16_inst_183_dout;
wire [8:8] rom16_inst_184_dout;
wire [9:9] rom16_inst_185_dout;
wire [10:10] rom16_inst_186_dout;
wire [11:11] rom16_inst_187_dout;
wire [12:12] rom16_inst_188_dout;
wire [13:13] rom16_inst_189_dout;
wire [14:14] rom16_inst_190_dout;
wire [15:15] rom16_inst_191_dout;
wire [0:0] rom16_inst_192_dout;
wire [1:1] rom16_inst_193_dout;
wire [2:2] rom16_inst_194_dout;
wire [3:3] rom16_inst_195_dout;
wire [4:4] rom16_inst_196_dout;
wire [5:5] rom16_inst_197_dout;
wire [6:6] rom16_inst_198_dout;
wire [7:7] rom16_inst_199_dout;
wire [8:8] rom16_inst_200_dout;
wire [9:9] rom16_inst_201_dout;
wire [10:10] rom16_inst_202_dout;
wire [11:11] rom16_inst_203_dout;
wire [12:12] rom16_inst_204_dout;
wire [13:13] rom16_inst_205_dout;
wire [14:14] rom16_inst_206_dout;
wire [15:15] rom16_inst_207_dout;
wire [0:0] rom16_inst_208_dout;
wire [1:1] rom16_inst_209_dout;
wire [2:2] rom16_inst_210_dout;
wire [3:3] rom16_inst_211_dout;
wire [4:4] rom16_inst_212_dout;
wire [5:5] rom16_inst_213_dout;
wire [6:6] rom16_inst_214_dout;
wire [7:7] rom16_inst_215_dout;
wire [8:8] rom16_inst_216_dout;
wire [9:9] rom16_inst_217_dout;
wire [10:10] rom16_inst_218_dout;
wire [11:11] rom16_inst_219_dout;
wire [12:12] rom16_inst_220_dout;
wire [13:13] rom16_inst_221_dout;
wire [14:14] rom16_inst_222_dout;
wire [15:15] rom16_inst_223_dout;
wire [0:0] rom16_inst_224_dout;
wire [1:1] rom16_inst_225_dout;
wire [2:2] rom16_inst_226_dout;
wire [3:3] rom16_inst_227_dout;
wire [4:4] rom16_inst_228_dout;
wire [5:5] rom16_inst_229_dout;
wire [6:6] rom16_inst_230_dout;
wire [7:7] rom16_inst_231_dout;
wire [8:8] rom16_inst_232_dout;
wire [9:9] rom16_inst_233_dout;
wire [10:10] rom16_inst_234_dout;
wire [11:11] rom16_inst_235_dout;
wire [12:12] rom16_inst_236_dout;
wire [13:13] rom16_inst_237_dout;
wire [14:14] rom16_inst_238_dout;
wire [15:15] rom16_inst_239_dout;
wire [0:0] rom16_inst_240_dout;
wire [1:1] rom16_inst_241_dout;
wire [2:2] rom16_inst_242_dout;
wire [3:3] rom16_inst_243_dout;
wire [4:4] rom16_inst_244_dout;
wire [5:5] rom16_inst_245_dout;
wire [6:6] rom16_inst_246_dout;
wire [7:7] rom16_inst_247_dout;
wire [8:8] rom16_inst_248_dout;
wire [9:9] rom16_inst_249_dout;
wire [10:10] rom16_inst_250_dout;
wire [11:11] rom16_inst_251_dout;
wire [12:12] rom16_inst_252_dout;
wire [13:13] rom16_inst_253_dout;
wire [14:14] rom16_inst_254_dout;
wire [15:15] rom16_inst_255_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_48;
wire mux_o_49;
wire mux_o_50;
wire mux_o_51;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_96;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_100;
wire mux_o_101;
wire mux_o_102;
wire mux_o_103;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_141;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_148;
wire mux_o_150;
wire mux_o_151;
wire mux_o_152;
wire mux_o_153;
wire mux_o_154;
wire mux_o_155;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_193;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_200;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_204;
wire mux_o_205;
wire mux_o_206;
wire mux_o_207;
wire mux_o_208;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;

ROM16 rom16_inst_0 (
    .DO(rom16_inst_0_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_0.INIT_0 = 16'h0000;

ROM16 rom16_inst_1 (
    .DO(rom16_inst_1_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_1.INIT_0 = 16'h0000;

ROM16 rom16_inst_2 (
    .DO(rom16_inst_2_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_2.INIT_0 = 16'h0000;

ROM16 rom16_inst_3 (
    .DO(rom16_inst_3_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_3.INIT_0 = 16'h0000;

ROM16 rom16_inst_4 (
    .DO(rom16_inst_4_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_4.INIT_0 = 16'h0000;

ROM16 rom16_inst_5 (
    .DO(rom16_inst_5_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_5.INIT_0 = 16'h6666;

ROM16 rom16_inst_6 (
    .DO(rom16_inst_6_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_6.INIT_0 = 16'hB4B4;

ROM16 rom16_inst_7 (
    .DO(rom16_inst_7_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_7.INIT_0 = 16'hC738;

ROM16 rom16_inst_8 (
    .DO(rom16_inst_8_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_8.INIT_0 = 16'h07C0;

ROM16 rom16_inst_9 (
    .DO(rom16_inst_9_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_9.INIT_0 = 16'hF800;

ROM16 rom16_inst_10 (
    .DO(rom16_inst_10_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_10.INIT_0 = 16'h0000;

ROM16 rom16_inst_11 (
    .DO(rom16_inst_11_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_11.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_12 (
    .DO(rom16_inst_12_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_12.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_13 (
    .DO(rom16_inst_13_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_13.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_14 (
    .DO(rom16_inst_14_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_14.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_15 (
    .DO(rom16_inst_15_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_15.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_16 (
    .DO(rom16_inst_16_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_16.INIT_0 = 16'h0000;

ROM16 rom16_inst_17 (
    .DO(rom16_inst_17_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_17.INIT_0 = 16'h0000;

ROM16 rom16_inst_18 (
    .DO(rom16_inst_18_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_18.INIT_0 = 16'h0000;

ROM16 rom16_inst_19 (
    .DO(rom16_inst_19_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_19.INIT_0 = 16'h0000;

ROM16 rom16_inst_20 (
    .DO(rom16_inst_20_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_20.INIT_0 = 16'h0000;

ROM16 rom16_inst_21 (
    .DO(rom16_inst_21_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_21.INIT_0 = 16'h6666;

ROM16 rom16_inst_22 (
    .DO(rom16_inst_22_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_22.INIT_0 = 16'hB4B4;

ROM16 rom16_inst_23 (
    .DO(rom16_inst_23_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_23.INIT_0 = 16'hC738;

ROM16 rom16_inst_24 (
    .DO(rom16_inst_24_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_24.INIT_0 = 16'hF83F;

ROM16 rom16_inst_25 (
    .DO(rom16_inst_25_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_25.INIT_0 = 16'h003F;

ROM16 rom16_inst_26 (
    .DO(rom16_inst_26_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_26.INIT_0 = 16'hFFC0;

ROM16 rom16_inst_27 (
    .DO(rom16_inst_27_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_27.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_28 (
    .DO(rom16_inst_28_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_28.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_29 (
    .DO(rom16_inst_29_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_29.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_30 (
    .DO(rom16_inst_30_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_30.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_31 (
    .DO(rom16_inst_31_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_31.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_32 (
    .DO(rom16_inst_32_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_32.INIT_0 = 16'h0000;

ROM16 rom16_inst_33 (
    .DO(rom16_inst_33_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_33.INIT_0 = 16'h0000;

ROM16 rom16_inst_34 (
    .DO(rom16_inst_34_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_34.INIT_0 = 16'h0000;

ROM16 rom16_inst_35 (
    .DO(rom16_inst_35_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_35.INIT_0 = 16'h0000;

ROM16 rom16_inst_36 (
    .DO(rom16_inst_36_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_36.INIT_0 = 16'h0000;

ROM16 rom16_inst_37 (
    .DO(rom16_inst_37_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_37.INIT_0 = 16'hFE66;

ROM16 rom16_inst_38 (
    .DO(rom16_inst_38_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_38.INIT_0 = 16'hFCB4;

ROM16 rom16_inst_39 (
    .DO(rom16_inst_39_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_39.INIT_0 = 16'hFF38;

ROM16 rom16_inst_40 (
    .DO(rom16_inst_40_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_40.INIT_0 = 16'hFFC0;

ROM16 rom16_inst_41 (
    .DO(rom16_inst_41_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_41.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_42 (
    .DO(rom16_inst_42_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_42.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_43 (
    .DO(rom16_inst_43_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_43.INIT_0 = 16'h4FFF;

ROM16 rom16_inst_44 (
    .DO(rom16_inst_44_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_44.INIT_0 = 16'h3FFF;

ROM16 rom16_inst_45 (
    .DO(rom16_inst_45_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_45.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_46 (
    .DO(rom16_inst_46_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_46.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_47 (
    .DO(rom16_inst_47_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_47.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_48 (
    .DO(rom16_inst_48_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_48.INIT_0 = 16'h0000;

ROM16 rom16_inst_49 (
    .DO(rom16_inst_49_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_49.INIT_0 = 16'h0000;

ROM16 rom16_inst_50 (
    .DO(rom16_inst_50_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_50.INIT_0 = 16'h0000;

ROM16 rom16_inst_51 (
    .DO(rom16_inst_51_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_51.INIT_0 = 16'h0000;

ROM16 rom16_inst_52 (
    .DO(rom16_inst_52_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_52.INIT_0 = 16'h0000;

ROM16 rom16_inst_53 (
    .DO(rom16_inst_53_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_53.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_54 (
    .DO(rom16_inst_54_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_54.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_55 (
    .DO(rom16_inst_55_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_55.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_56 (
    .DO(rom16_inst_56_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_56.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_57 (
    .DO(rom16_inst_57_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_57.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_58 (
    .DO(rom16_inst_58_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_58.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_59 (
    .DO(rom16_inst_59_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_59.INIT_0 = 16'h4B4B;

ROM16 rom16_inst_60 (
    .DO(rom16_inst_60_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_60.INIT_0 = 16'h38C7;

ROM16 rom16_inst_61 (
    .DO(rom16_inst_61_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_61.INIT_0 = 16'h07C0;

ROM16 rom16_inst_62 (
    .DO(rom16_inst_62_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_62.INIT_0 = 16'h003F;

ROM16 rom16_inst_63 (
    .DO(rom16_inst_63_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_63.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_64 (
    .DO(rom16_inst_64_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_64.INIT_0 = 16'h0000;

ROM16 rom16_inst_65 (
    .DO(rom16_inst_65_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_65.INIT_0 = 16'h0000;

ROM16 rom16_inst_66 (
    .DO(rom16_inst_66_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_66.INIT_0 = 16'h0000;

ROM16 rom16_inst_67 (
    .DO(rom16_inst_67_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_67.INIT_0 = 16'h0000;

ROM16 rom16_inst_68 (
    .DO(rom16_inst_68_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_68.INIT_0 = 16'h0000;

ROM16 rom16_inst_69 (
    .DO(rom16_inst_69_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_69.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_70 (
    .DO(rom16_inst_70_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_70.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_71 (
    .DO(rom16_inst_71_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_71.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_72 (
    .DO(rom16_inst_72_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_72.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_73 (
    .DO(rom16_inst_73_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_73.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_74 (
    .DO(rom16_inst_74_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_74.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_75 (
    .DO(rom16_inst_75_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_75.INIT_0 = 16'h4B4B;

ROM16 rom16_inst_76 (
    .DO(rom16_inst_76_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_76.INIT_0 = 16'h38C7;

ROM16 rom16_inst_77 (
    .DO(rom16_inst_77_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_77.INIT_0 = 16'hF83F;

ROM16 rom16_inst_78 (
    .DO(rom16_inst_78_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_78.INIT_0 = 16'h07FF;

ROM16 rom16_inst_79 (
    .DO(rom16_inst_79_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_79.INIT_0 = 16'h0000;

ROM16 rom16_inst_80 (
    .DO(rom16_inst_80_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_80.INIT_0 = 16'h9680;

ROM16 rom16_inst_81 (
    .DO(rom16_inst_81_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_81.INIT_0 = 16'hE700;

ROM16 rom16_inst_82 (
    .DO(rom16_inst_82_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_82.INIT_0 = 16'hF800;

ROM16 rom16_inst_83 (
    .DO(rom16_inst_83_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_83.INIT_0 = 16'h0000;

ROM16 rom16_inst_84 (
    .DO(rom16_inst_84_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_84.INIT_0 = 16'h0000;

ROM16 rom16_inst_85 (
    .DO(rom16_inst_85_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_85.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_86 (
    .DO(rom16_inst_86_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_86.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_87 (
    .DO(rom16_inst_87_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_87.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_88 (
    .DO(rom16_inst_88_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_88.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_89 (
    .DO(rom16_inst_89_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_89.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_90 (
    .DO(rom16_inst_90_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_90.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_91 (
    .DO(rom16_inst_91_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_91.INIT_0 = 16'h000B;

ROM16 rom16_inst_92 (
    .DO(rom16_inst_92_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_92.INIT_0 = 16'h0007;

ROM16 rom16_inst_93 (
    .DO(rom16_inst_93_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_93.INIT_0 = 16'h0000;

ROM16 rom16_inst_94 (
    .DO(rom16_inst_94_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_94.INIT_0 = 16'h0000;

ROM16 rom16_inst_95 (
    .DO(rom16_inst_95_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_95.INIT_0 = 16'h0000;

ROM16 rom16_inst_96 (
    .DO(rom16_inst_96_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_96.INIT_0 = 16'h9696;

ROM16 rom16_inst_97 (
    .DO(rom16_inst_97_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_97.INIT_0 = 16'hE718;

ROM16 rom16_inst_98 (
    .DO(rom16_inst_98_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_98.INIT_0 = 16'h07E0;

ROM16 rom16_inst_99 (
    .DO(rom16_inst_99_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_99.INIT_0 = 16'h07FF;

ROM16 rom16_inst_100 (
    .DO(rom16_inst_100_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_100.INIT_0 = 16'hF800;

ROM16 rom16_inst_101 (
    .DO(rom16_inst_101_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_101.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_102 (
    .DO(rom16_inst_102_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_102.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_103 (
    .DO(rom16_inst_103_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_103.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_104 (
    .DO(rom16_inst_104_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_104.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_105 (
    .DO(rom16_inst_105_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_105.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_106 (
    .DO(rom16_inst_106_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_106.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_107 (
    .DO(rom16_inst_107_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_107.INIT_0 = 16'h0000;

ROM16 rom16_inst_108 (
    .DO(rom16_inst_108_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_108.INIT_0 = 16'h0000;

ROM16 rom16_inst_109 (
    .DO(rom16_inst_109_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_109.INIT_0 = 16'h0000;

ROM16 rom16_inst_110 (
    .DO(rom16_inst_110_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_110.INIT_0 = 16'h0000;

ROM16 rom16_inst_111 (
    .DO(rom16_inst_111_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_111.INIT_0 = 16'h0000;

ROM16 rom16_inst_112 (
    .DO(rom16_inst_112_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_112.INIT_0 = 16'h9696;

ROM16 rom16_inst_113 (
    .DO(rom16_inst_113_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_113.INIT_0 = 16'hE718;

ROM16 rom16_inst_114 (
    .DO(rom16_inst_114_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_114.INIT_0 = 16'hF81F;

ROM16 rom16_inst_115 (
    .DO(rom16_inst_115_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_115.INIT_0 = 16'hFFE0;

ROM16 rom16_inst_116 (
    .DO(rom16_inst_116_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_116.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_117 (
    .DO(rom16_inst_117_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_117.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_118 (
    .DO(rom16_inst_118_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_118.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_119 (
    .DO(rom16_inst_119_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_119.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_120 (
    .DO(rom16_inst_120_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_120.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_121 (
    .DO(rom16_inst_121_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_121.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_122 (
    .DO(rom16_inst_122_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_122.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_123 (
    .DO(rom16_inst_123_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_123.INIT_0 = 16'h0000;

ROM16 rom16_inst_124 (
    .DO(rom16_inst_124_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_124.INIT_0 = 16'h0000;

ROM16 rom16_inst_125 (
    .DO(rom16_inst_125_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_125.INIT_0 = 16'h0000;

ROM16 rom16_inst_126 (
    .DO(rom16_inst_126_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_126.INIT_0 = 16'h0000;

ROM16 rom16_inst_127 (
    .DO(rom16_inst_127_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_127.INIT_0 = 16'h0000;

ROM16 rom16_inst_128 (
    .DO(rom16_inst_128_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_128.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_129 (
    .DO(rom16_inst_129_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_129.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_130 (
    .DO(rom16_inst_130_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_130.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_131 (
    .DO(rom16_inst_131_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_131.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_132 (
    .DO(rom16_inst_132_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_132.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_133 (
    .DO(rom16_inst_133_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_133.INIT_0 = 16'h3333;

ROM16 rom16_inst_134 (
    .DO(rom16_inst_134_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_134.INIT_0 = 16'h6969;

ROM16 rom16_inst_135 (
    .DO(rom16_inst_135_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_135.INIT_0 = 16'h18E7;

ROM16 rom16_inst_136 (
    .DO(rom16_inst_136_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_136.INIT_0 = 16'hF81F;

ROM16 rom16_inst_137 (
    .DO(rom16_inst_137_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_137.INIT_0 = 16'h07FF;

ROM16 rom16_inst_138 (
    .DO(rom16_inst_138_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_138.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_139 (
    .DO(rom16_inst_139_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_139.INIT_0 = 16'h0000;

ROM16 rom16_inst_140 (
    .DO(rom16_inst_140_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_140.INIT_0 = 16'h0000;

ROM16 rom16_inst_141 (
    .DO(rom16_inst_141_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_141.INIT_0 = 16'h0000;

ROM16 rom16_inst_142 (
    .DO(rom16_inst_142_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_142.INIT_0 = 16'h0000;

ROM16 rom16_inst_143 (
    .DO(rom16_inst_143_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_143.INIT_0 = 16'h0000;

ROM16 rom16_inst_144 (
    .DO(rom16_inst_144_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_144.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_145 (
    .DO(rom16_inst_145_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_145.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_146 (
    .DO(rom16_inst_146_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_146.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_147 (
    .DO(rom16_inst_147_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_147.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_148 (
    .DO(rom16_inst_148_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_148.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_149 (
    .DO(rom16_inst_149_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_149.INIT_0 = 16'h3333;

ROM16 rom16_inst_150 (
    .DO(rom16_inst_150_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_150.INIT_0 = 16'h6969;

ROM16 rom16_inst_151 (
    .DO(rom16_inst_151_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_151.INIT_0 = 16'h18E7;

ROM16 rom16_inst_152 (
    .DO(rom16_inst_152_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_152.INIT_0 = 16'h07E0;

ROM16 rom16_inst_153 (
    .DO(rom16_inst_153_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_153.INIT_0 = 16'hFFE0;

ROM16 rom16_inst_154 (
    .DO(rom16_inst_154_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_154.INIT_0 = 16'h001F;

ROM16 rom16_inst_155 (
    .DO(rom16_inst_155_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_155.INIT_0 = 16'h0000;

ROM16 rom16_inst_156 (
    .DO(rom16_inst_156_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_156.INIT_0 = 16'h0000;

ROM16 rom16_inst_157 (
    .DO(rom16_inst_157_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_157.INIT_0 = 16'h0000;

ROM16 rom16_inst_158 (
    .DO(rom16_inst_158_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_158.INIT_0 = 16'h0000;

ROM16 rom16_inst_159 (
    .DO(rom16_inst_159_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_159.INIT_0 = 16'h0000;

ROM16 rom16_inst_160 (
    .DO(rom16_inst_160_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_160.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_161 (
    .DO(rom16_inst_161_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_161.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_162 (
    .DO(rom16_inst_162_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_162.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_163 (
    .DO(rom16_inst_163_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_163.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_164 (
    .DO(rom16_inst_164_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_164.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_165 (
    .DO(rom16_inst_165_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_165.INIT_0 = 16'h0333;

ROM16 rom16_inst_166 (
    .DO(rom16_inst_166_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_166.INIT_0 = 16'h0169;

ROM16 rom16_inst_167 (
    .DO(rom16_inst_167_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_167.INIT_0 = 16'h00E7;

ROM16 rom16_inst_168 (
    .DO(rom16_inst_168_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_168.INIT_0 = 16'h001F;

ROM16 rom16_inst_169 (
    .DO(rom16_inst_169_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_169.INIT_0 = 16'h0000;

ROM16 rom16_inst_170 (
    .DO(rom16_inst_170_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_170.INIT_0 = 16'h0000;

ROM16 rom16_inst_171 (
    .DO(rom16_inst_171_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_171.INIT_0 = 16'hD000;

ROM16 rom16_inst_172 (
    .DO(rom16_inst_172_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_172.INIT_0 = 16'hE000;

ROM16 rom16_inst_173 (
    .DO(rom16_inst_173_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_173.INIT_0 = 16'h0000;

ROM16 rom16_inst_174 (
    .DO(rom16_inst_174_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_174.INIT_0 = 16'h0000;

ROM16 rom16_inst_175 (
    .DO(rom16_inst_175_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_175.INIT_0 = 16'h0000;

ROM16 rom16_inst_176 (
    .DO(rom16_inst_176_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_176.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_177 (
    .DO(rom16_inst_177_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_177.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_178 (
    .DO(rom16_inst_178_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_178.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_179 (
    .DO(rom16_inst_179_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_179.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_180 (
    .DO(rom16_inst_180_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_180.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_181 (
    .DO(rom16_inst_181_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_181.INIT_0 = 16'h0000;

ROM16 rom16_inst_182 (
    .DO(rom16_inst_182_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_182.INIT_0 = 16'h0000;

ROM16 rom16_inst_183 (
    .DO(rom16_inst_183_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_183.INIT_0 = 16'h0000;

ROM16 rom16_inst_184 (
    .DO(rom16_inst_184_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_184.INIT_0 = 16'h0000;

ROM16 rom16_inst_185 (
    .DO(rom16_inst_185_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_185.INIT_0 = 16'h0000;

ROM16 rom16_inst_186 (
    .DO(rom16_inst_186_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_186.INIT_0 = 16'h0000;

ROM16 rom16_inst_187 (
    .DO(rom16_inst_187_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_187.INIT_0 = 16'hD2D2;

ROM16 rom16_inst_188 (
    .DO(rom16_inst_188_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_188.INIT_0 = 16'hE31C;

ROM16 rom16_inst_189 (
    .DO(rom16_inst_189_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_189.INIT_0 = 16'hFC1F;

ROM16 rom16_inst_190 (
    .DO(rom16_inst_190_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_190.INIT_0 = 16'hFFE0;

ROM16 rom16_inst_191 (
    .DO(rom16_inst_191_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_191.INIT_0 = 16'h0000;

ROM16 rom16_inst_192 (
    .DO(rom16_inst_192_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_192.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_193 (
    .DO(rom16_inst_193_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_193.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_194 (
    .DO(rom16_inst_194_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_194.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_195 (
    .DO(rom16_inst_195_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_195.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_196 (
    .DO(rom16_inst_196_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_196.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_197 (
    .DO(rom16_inst_197_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_197.INIT_0 = 16'h0000;

ROM16 rom16_inst_198 (
    .DO(rom16_inst_198_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_198.INIT_0 = 16'h0000;

ROM16 rom16_inst_199 (
    .DO(rom16_inst_199_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_199.INIT_0 = 16'h0000;

ROM16 rom16_inst_200 (
    .DO(rom16_inst_200_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_200.INIT_0 = 16'h0000;

ROM16 rom16_inst_201 (
    .DO(rom16_inst_201_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_201.INIT_0 = 16'h0000;

ROM16 rom16_inst_202 (
    .DO(rom16_inst_202_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_202.INIT_0 = 16'h0000;

ROM16 rom16_inst_203 (
    .DO(rom16_inst_203_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_203.INIT_0 = 16'hD2D2;

ROM16 rom16_inst_204 (
    .DO(rom16_inst_204_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_204.INIT_0 = 16'hE31C;

ROM16 rom16_inst_205 (
    .DO(rom16_inst_205_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_205.INIT_0 = 16'h03E0;

ROM16 rom16_inst_206 (
    .DO(rom16_inst_206_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_206.INIT_0 = 16'hFC00;

ROM16 rom16_inst_207 (
    .DO(rom16_inst_207_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_207.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_208 (
    .DO(rom16_inst_208_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_208.INIT_0 = 16'h2D3F;

ROM16 rom16_inst_209 (
    .DO(rom16_inst_209_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_209.INIT_0 = 16'h1CFF;

ROM16 rom16_inst_210 (
    .DO(rom16_inst_210_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_210.INIT_0 = 16'h03FF;

ROM16 rom16_inst_211 (
    .DO(rom16_inst_211_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_211.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_212 (
    .DO(rom16_inst_212_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_212.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_213 (
    .DO(rom16_inst_213_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_213.INIT_0 = 16'h0000;

ROM16 rom16_inst_214 (
    .DO(rom16_inst_214_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_214.INIT_0 = 16'h0000;

ROM16 rom16_inst_215 (
    .DO(rom16_inst_215_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_215.INIT_0 = 16'h0000;

ROM16 rom16_inst_216 (
    .DO(rom16_inst_216_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_216.INIT_0 = 16'h0000;

ROM16 rom16_inst_217 (
    .DO(rom16_inst_217_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_217.INIT_0 = 16'h0000;

ROM16 rom16_inst_218 (
    .DO(rom16_inst_218_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_218.INIT_0 = 16'h0000;

ROM16 rom16_inst_219 (
    .DO(rom16_inst_219_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_219.INIT_0 = 16'hFFF2;

ROM16 rom16_inst_220 (
    .DO(rom16_inst_220_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_220.INIT_0 = 16'hFFFC;

ROM16 rom16_inst_221 (
    .DO(rom16_inst_221_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_221.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_222 (
    .DO(rom16_inst_222_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_222.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_223 (
    .DO(rom16_inst_223_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_223.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_224 (
    .DO(rom16_inst_224_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_224.INIT_0 = 16'h2D2D;

ROM16 rom16_inst_225 (
    .DO(rom16_inst_225_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_225.INIT_0 = 16'h1CE3;

ROM16 rom16_inst_226 (
    .DO(rom16_inst_226_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_226.INIT_0 = 16'hFC1F;

ROM16 rom16_inst_227 (
    .DO(rom16_inst_227_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_227.INIT_0 = 16'hFC00;

ROM16 rom16_inst_228 (
    .DO(rom16_inst_228_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_228.INIT_0 = 16'h03FF;

ROM16 rom16_inst_229 (
    .DO(rom16_inst_229_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_229.INIT_0 = 16'h0000;

ROM16 rom16_inst_230 (
    .DO(rom16_inst_230_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_230.INIT_0 = 16'h0000;

ROM16 rom16_inst_231 (
    .DO(rom16_inst_231_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_231.INIT_0 = 16'h0000;

ROM16 rom16_inst_232 (
    .DO(rom16_inst_232_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_232.INIT_0 = 16'h0000;

ROM16 rom16_inst_233 (
    .DO(rom16_inst_233_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_233.INIT_0 = 16'h0000;

ROM16 rom16_inst_234 (
    .DO(rom16_inst_234_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_234.INIT_0 = 16'h0000;

ROM16 rom16_inst_235 (
    .DO(rom16_inst_235_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_235.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_236 (
    .DO(rom16_inst_236_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_236.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_237 (
    .DO(rom16_inst_237_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_237.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_238 (
    .DO(rom16_inst_238_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_238.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_239 (
    .DO(rom16_inst_239_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_239.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_240 (
    .DO(rom16_inst_240_dout[0]),
    .AD(ad[3:0])
);

defparam rom16_inst_240.INIT_0 = 16'h2D2D;

ROM16 rom16_inst_241 (
    .DO(rom16_inst_241_dout[1]),
    .AD(ad[3:0])
);

defparam rom16_inst_241.INIT_0 = 16'h1CE3;

ROM16 rom16_inst_242 (
    .DO(rom16_inst_242_dout[2]),
    .AD(ad[3:0])
);

defparam rom16_inst_242.INIT_0 = 16'h03E0;

ROM16 rom16_inst_243 (
    .DO(rom16_inst_243_dout[3]),
    .AD(ad[3:0])
);

defparam rom16_inst_243.INIT_0 = 16'h001F;

ROM16 rom16_inst_244 (
    .DO(rom16_inst_244_dout[4]),
    .AD(ad[3:0])
);

defparam rom16_inst_244.INIT_0 = 16'h0000;

ROM16 rom16_inst_245 (
    .DO(rom16_inst_245_dout[5]),
    .AD(ad[3:0])
);

defparam rom16_inst_245.INIT_0 = 16'h0000;

ROM16 rom16_inst_246 (
    .DO(rom16_inst_246_dout[6]),
    .AD(ad[3:0])
);

defparam rom16_inst_246.INIT_0 = 16'h0000;

ROM16 rom16_inst_247 (
    .DO(rom16_inst_247_dout[7]),
    .AD(ad[3:0])
);

defparam rom16_inst_247.INIT_0 = 16'h0000;

ROM16 rom16_inst_248 (
    .DO(rom16_inst_248_dout[8]),
    .AD(ad[3:0])
);

defparam rom16_inst_248.INIT_0 = 16'h0000;

ROM16 rom16_inst_249 (
    .DO(rom16_inst_249_dout[9]),
    .AD(ad[3:0])
);

defparam rom16_inst_249.INIT_0 = 16'h0000;

ROM16 rom16_inst_250 (
    .DO(rom16_inst_250_dout[10]),
    .AD(ad[3:0])
);

defparam rom16_inst_250.INIT_0 = 16'h0000;

ROM16 rom16_inst_251 (
    .DO(rom16_inst_251_dout[11]),
    .AD(ad[3:0])
);

defparam rom16_inst_251.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_252 (
    .DO(rom16_inst_252_dout[12]),
    .AD(ad[3:0])
);

defparam rom16_inst_252.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_253 (
    .DO(rom16_inst_253_dout[13]),
    .AD(ad[3:0])
);

defparam rom16_inst_253.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_254 (
    .DO(rom16_inst_254_dout[14]),
    .AD(ad[3:0])
);

defparam rom16_inst_254.INIT_0 = 16'hFFFF;

ROM16 rom16_inst_255 (
    .DO(rom16_inst_255_dout[15]),
    .AD(ad[3:0])
);

defparam rom16_inst_255.INIT_0 = 16'hFFFF;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(rom16_inst_0_dout[0]),
  .I1(rom16_inst_16_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(rom16_inst_32_dout[0]),
  .I1(rom16_inst_48_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(rom16_inst_64_dout[0]),
  .I1(rom16_inst_80_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(rom16_inst_96_dout[0]),
  .I1(rom16_inst_112_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(rom16_inst_128_dout[0]),
  .I1(rom16_inst_144_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(rom16_inst_160_dout[0]),
  .I1(rom16_inst_176_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(rom16_inst_192_dout[0]),
  .I1(rom16_inst_208_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(rom16_inst_224_dout[0]),
  .I1(rom16_inst_240_dout[0]),
  .S0(ad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(ad[5])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(ad[5])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(ad[5])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(ad[5])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(ad[6])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(ad[6])
);
MUX2 mux_inst_14 (
  .O(dout[0]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(ad[7])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(rom16_inst_1_dout[1]),
  .I1(rom16_inst_17_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(rom16_inst_33_dout[1]),
  .I1(rom16_inst_49_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(rom16_inst_65_dout[1]),
  .I1(rom16_inst_81_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(rom16_inst_97_dout[1]),
  .I1(rom16_inst_113_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(rom16_inst_129_dout[1]),
  .I1(rom16_inst_145_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(rom16_inst_161_dout[1]),
  .I1(rom16_inst_177_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(rom16_inst_193_dout[1]),
  .I1(rom16_inst_209_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(rom16_inst_225_dout[1]),
  .I1(rom16_inst_241_dout[1]),
  .S0(ad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(ad[5])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(mux_o_17),
  .I1(mux_o_18),
  .S0(ad[5])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_19),
  .I1(mux_o_20),
  .S0(ad[5])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(ad[5])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_23),
  .I1(mux_o_24),
  .S0(ad[6])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(ad[6])
);
MUX2 mux_inst_29 (
  .O(dout[1]),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(ad[7])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(rom16_inst_2_dout[2]),
  .I1(rom16_inst_18_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(rom16_inst_34_dout[2]),
  .I1(rom16_inst_50_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(rom16_inst_66_dout[2]),
  .I1(rom16_inst_82_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(rom16_inst_98_dout[2]),
  .I1(rom16_inst_114_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(rom16_inst_130_dout[2]),
  .I1(rom16_inst_146_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(rom16_inst_162_dout[2]),
  .I1(rom16_inst_178_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(rom16_inst_194_dout[2]),
  .I1(rom16_inst_210_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(rom16_inst_226_dout[2]),
  .I1(rom16_inst_242_dout[2]),
  .S0(ad[4])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_30),
  .I1(mux_o_31),
  .S0(ad[5])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_32),
  .I1(mux_o_33),
  .S0(ad[5])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_34),
  .I1(mux_o_35),
  .S0(ad[5])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(ad[5])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(ad[6])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(ad[6])
);
MUX2 mux_inst_44 (
  .O(dout[2]),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(ad[7])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(rom16_inst_3_dout[3]),
  .I1(rom16_inst_19_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(rom16_inst_35_dout[3]),
  .I1(rom16_inst_51_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(rom16_inst_67_dout[3]),
  .I1(rom16_inst_83_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_48 (
  .O(mux_o_48),
  .I0(rom16_inst_99_dout[3]),
  .I1(rom16_inst_115_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(rom16_inst_131_dout[3]),
  .I1(rom16_inst_147_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(rom16_inst_163_dout[3]),
  .I1(rom16_inst_179_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_51 (
  .O(mux_o_51),
  .I0(rom16_inst_195_dout[3]),
  .I1(rom16_inst_211_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(rom16_inst_227_dout[3]),
  .I1(rom16_inst_243_dout[3]),
  .S0(ad[4])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(ad[5])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(mux_o_47),
  .I1(mux_o_48),
  .S0(ad[5])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(ad[5])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(mux_o_51),
  .I1(mux_o_52),
  .S0(ad[5])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(mux_o_53),
  .I1(mux_o_54),
  .S0(ad[6])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(mux_o_55),
  .I1(mux_o_56),
  .S0(ad[6])
);
MUX2 mux_inst_59 (
  .O(dout[3]),
  .I0(mux_o_57),
  .I1(mux_o_58),
  .S0(ad[7])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(rom16_inst_4_dout[4]),
  .I1(rom16_inst_20_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(rom16_inst_36_dout[4]),
  .I1(rom16_inst_52_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(rom16_inst_68_dout[4]),
  .I1(rom16_inst_84_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(rom16_inst_100_dout[4]),
  .I1(rom16_inst_116_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(rom16_inst_132_dout[4]),
  .I1(rom16_inst_148_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(rom16_inst_164_dout[4]),
  .I1(rom16_inst_180_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(rom16_inst_196_dout[4]),
  .I1(rom16_inst_212_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(rom16_inst_228_dout[4]),
  .I1(rom16_inst_244_dout[4]),
  .S0(ad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(ad[5])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(ad[5])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(ad[5])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(ad[5])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(ad[6])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(ad[6])
);
MUX2 mux_inst_74 (
  .O(dout[4]),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(ad[7])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(rom16_inst_5_dout[5]),
  .I1(rom16_inst_21_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(rom16_inst_37_dout[5]),
  .I1(rom16_inst_53_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(rom16_inst_69_dout[5]),
  .I1(rom16_inst_85_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(rom16_inst_101_dout[5]),
  .I1(rom16_inst_117_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(rom16_inst_133_dout[5]),
  .I1(rom16_inst_149_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(rom16_inst_165_dout[5]),
  .I1(rom16_inst_181_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(rom16_inst_197_dout[5]),
  .I1(rom16_inst_213_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(rom16_inst_229_dout[5]),
  .I1(rom16_inst_245_dout[5]),
  .S0(ad[4])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_75),
  .I1(mux_o_76),
  .S0(ad[5])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(ad[5])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(ad[5])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(ad[5])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(ad[6])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(ad[6])
);
MUX2 mux_inst_89 (
  .O(dout[5]),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(ad[7])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(rom16_inst_6_dout[6]),
  .I1(rom16_inst_22_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(rom16_inst_38_dout[6]),
  .I1(rom16_inst_54_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(rom16_inst_70_dout[6]),
  .I1(rom16_inst_86_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(rom16_inst_102_dout[6]),
  .I1(rom16_inst_118_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(rom16_inst_134_dout[6]),
  .I1(rom16_inst_150_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(rom16_inst_166_dout[6]),
  .I1(rom16_inst_182_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_96 (
  .O(mux_o_96),
  .I0(rom16_inst_198_dout[6]),
  .I1(rom16_inst_214_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(rom16_inst_230_dout[6]),
  .I1(rom16_inst_246_dout[6]),
  .S0(ad[4])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(ad[5])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(ad[5])
);
MUX2 mux_inst_100 (
  .O(mux_o_100),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(ad[5])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_96),
  .I1(mux_o_97),
  .S0(ad[5])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_98),
  .I1(mux_o_99),
  .S0(ad[6])
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(mux_o_100),
  .I1(mux_o_101),
  .S0(ad[6])
);
MUX2 mux_inst_104 (
  .O(dout[6]),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(ad[7])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(rom16_inst_7_dout[7]),
  .I1(rom16_inst_23_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(rom16_inst_39_dout[7]),
  .I1(rom16_inst_55_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(rom16_inst_71_dout[7]),
  .I1(rom16_inst_87_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(rom16_inst_103_dout[7]),
  .I1(rom16_inst_119_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(rom16_inst_135_dout[7]),
  .I1(rom16_inst_151_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(rom16_inst_167_dout[7]),
  .I1(rom16_inst_183_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(rom16_inst_199_dout[7]),
  .I1(rom16_inst_215_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(rom16_inst_231_dout[7]),
  .I1(rom16_inst_247_dout[7]),
  .S0(ad[4])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(mux_o_105),
  .I1(mux_o_106),
  .S0(ad[5])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(mux_o_107),
  .I1(mux_o_108),
  .S0(ad[5])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(mux_o_109),
  .I1(mux_o_110),
  .S0(ad[5])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(mux_o_111),
  .I1(mux_o_112),
  .S0(ad[5])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(mux_o_113),
  .I1(mux_o_114),
  .S0(ad[6])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(mux_o_115),
  .I1(mux_o_116),
  .S0(ad[6])
);
MUX2 mux_inst_119 (
  .O(dout[7]),
  .I0(mux_o_117),
  .I1(mux_o_118),
  .S0(ad[7])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(rom16_inst_8_dout[8]),
  .I1(rom16_inst_24_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(rom16_inst_40_dout[8]),
  .I1(rom16_inst_56_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(rom16_inst_72_dout[8]),
  .I1(rom16_inst_88_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(rom16_inst_104_dout[8]),
  .I1(rom16_inst_120_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(rom16_inst_136_dout[8]),
  .I1(rom16_inst_152_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(rom16_inst_168_dout[8]),
  .I1(rom16_inst_184_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(rom16_inst_200_dout[8]),
  .I1(rom16_inst_216_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(rom16_inst_232_dout[8]),
  .I1(rom16_inst_248_dout[8]),
  .S0(ad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(ad[5])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(ad[5])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(ad[5])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(ad[5])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_128),
  .I1(mux_o_129),
  .S0(ad[6])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_130),
  .I1(mux_o_131),
  .S0(ad[6])
);
MUX2 mux_inst_134 (
  .O(dout[8]),
  .I0(mux_o_132),
  .I1(mux_o_133),
  .S0(ad[7])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(rom16_inst_9_dout[9]),
  .I1(rom16_inst_25_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(rom16_inst_41_dout[9]),
  .I1(rom16_inst_57_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(rom16_inst_73_dout[9]),
  .I1(rom16_inst_89_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(rom16_inst_105_dout[9]),
  .I1(rom16_inst_121_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(rom16_inst_137_dout[9]),
  .I1(rom16_inst_153_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(rom16_inst_169_dout[9]),
  .I1(rom16_inst_185_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_141 (
  .O(mux_o_141),
  .I0(rom16_inst_201_dout[9]),
  .I1(rom16_inst_217_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(rom16_inst_233_dout[9]),
  .I1(rom16_inst_249_dout[9]),
  .S0(ad[4])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(ad[5])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(ad[5])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(ad[5])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_141),
  .I1(mux_o_142),
  .S0(ad[5])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_143),
  .I1(mux_o_144),
  .S0(ad[6])
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(mux_o_145),
  .I1(mux_o_146),
  .S0(ad[6])
);
MUX2 mux_inst_149 (
  .O(dout[9]),
  .I0(mux_o_147),
  .I1(mux_o_148),
  .S0(ad[7])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(rom16_inst_10_dout[10]),
  .I1(rom16_inst_26_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(rom16_inst_42_dout[10]),
  .I1(rom16_inst_58_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_152 (
  .O(mux_o_152),
  .I0(rom16_inst_74_dout[10]),
  .I1(rom16_inst_90_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(rom16_inst_106_dout[10]),
  .I1(rom16_inst_122_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(rom16_inst_138_dout[10]),
  .I1(rom16_inst_154_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(rom16_inst_170_dout[10]),
  .I1(rom16_inst_186_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(rom16_inst_202_dout[10]),
  .I1(rom16_inst_218_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(rom16_inst_234_dout[10]),
  .I1(rom16_inst_250_dout[10]),
  .S0(ad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(ad[5])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(mux_o_152),
  .I1(mux_o_153),
  .S0(ad[5])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(ad[5])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(ad[5])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(ad[6])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(ad[6])
);
MUX2 mux_inst_164 (
  .O(dout[10]),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(ad[7])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(rom16_inst_11_dout[11]),
  .I1(rom16_inst_27_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(rom16_inst_43_dout[11]),
  .I1(rom16_inst_59_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(rom16_inst_75_dout[11]),
  .I1(rom16_inst_91_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(rom16_inst_107_dout[11]),
  .I1(rom16_inst_123_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(rom16_inst_139_dout[11]),
  .I1(rom16_inst_155_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(rom16_inst_171_dout[11]),
  .I1(rom16_inst_187_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(rom16_inst_203_dout[11]),
  .I1(rom16_inst_219_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(rom16_inst_235_dout[11]),
  .I1(rom16_inst_251_dout[11]),
  .S0(ad[4])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(mux_o_165),
  .I1(mux_o_166),
  .S0(ad[5])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(mux_o_167),
  .I1(mux_o_168),
  .S0(ad[5])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(mux_o_169),
  .I1(mux_o_170),
  .S0(ad[5])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(ad[5])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(ad[6])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_175),
  .I1(mux_o_176),
  .S0(ad[6])
);
MUX2 mux_inst_179 (
  .O(dout[11]),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(ad[7])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(rom16_inst_12_dout[12]),
  .I1(rom16_inst_28_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(rom16_inst_44_dout[12]),
  .I1(rom16_inst_60_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(rom16_inst_76_dout[12]),
  .I1(rom16_inst_92_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(rom16_inst_108_dout[12]),
  .I1(rom16_inst_124_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(rom16_inst_140_dout[12]),
  .I1(rom16_inst_156_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(rom16_inst_172_dout[12]),
  .I1(rom16_inst_188_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(rom16_inst_204_dout[12]),
  .I1(rom16_inst_220_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(rom16_inst_236_dout[12]),
  .I1(rom16_inst_252_dout[12]),
  .S0(ad[4])
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(mux_o_180),
  .I1(mux_o_181),
  .S0(ad[5])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_182),
  .I1(mux_o_183),
  .S0(ad[5])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_184),
  .I1(mux_o_185),
  .S0(ad[5])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_186),
  .I1(mux_o_187),
  .S0(ad[5])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_188),
  .I1(mux_o_189),
  .S0(ad[6])
);
MUX2 mux_inst_193 (
  .O(mux_o_193),
  .I0(mux_o_190),
  .I1(mux_o_191),
  .S0(ad[6])
);
MUX2 mux_inst_194 (
  .O(dout[12]),
  .I0(mux_o_192),
  .I1(mux_o_193),
  .S0(ad[7])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(rom16_inst_13_dout[13]),
  .I1(rom16_inst_29_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(rom16_inst_45_dout[13]),
  .I1(rom16_inst_61_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(rom16_inst_77_dout[13]),
  .I1(rom16_inst_93_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(rom16_inst_109_dout[13]),
  .I1(rom16_inst_125_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(rom16_inst_141_dout[13]),
  .I1(rom16_inst_157_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(rom16_inst_173_dout[13]),
  .I1(rom16_inst_189_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(rom16_inst_205_dout[13]),
  .I1(rom16_inst_221_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(rom16_inst_237_dout[13]),
  .I1(rom16_inst_253_dout[13]),
  .S0(ad[4])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_195),
  .I1(mux_o_196),
  .S0(ad[5])
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_197),
  .I1(mux_o_198),
  .S0(ad[5])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_199),
  .I1(mux_o_200),
  .S0(ad[5])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(ad[5])
);
MUX2 mux_inst_207 (
  .O(mux_o_207),
  .I0(mux_o_203),
  .I1(mux_o_204),
  .S0(ad[6])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(ad[6])
);
MUX2 mux_inst_209 (
  .O(dout[13]),
  .I0(mux_o_207),
  .I1(mux_o_208),
  .S0(ad[7])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(rom16_inst_14_dout[14]),
  .I1(rom16_inst_30_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(rom16_inst_46_dout[14]),
  .I1(rom16_inst_62_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(rom16_inst_78_dout[14]),
  .I1(rom16_inst_94_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(rom16_inst_110_dout[14]),
  .I1(rom16_inst_126_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(rom16_inst_142_dout[14]),
  .I1(rom16_inst_158_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(rom16_inst_174_dout[14]),
  .I1(rom16_inst_190_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(rom16_inst_206_dout[14]),
  .I1(rom16_inst_222_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(rom16_inst_238_dout[14]),
  .I1(rom16_inst_254_dout[14]),
  .S0(ad[4])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(ad[5])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(ad[5])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(ad[5])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(ad[5])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(ad[6])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(ad[6])
);
MUX2 mux_inst_224 (
  .O(dout[14]),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(ad[7])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(rom16_inst_15_dout[15]),
  .I1(rom16_inst_31_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(rom16_inst_47_dout[15]),
  .I1(rom16_inst_63_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(rom16_inst_79_dout[15]),
  .I1(rom16_inst_95_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(rom16_inst_111_dout[15]),
  .I1(rom16_inst_127_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(rom16_inst_143_dout[15]),
  .I1(rom16_inst_159_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(rom16_inst_175_dout[15]),
  .I1(rom16_inst_191_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(rom16_inst_207_dout[15]),
  .I1(rom16_inst_223_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(rom16_inst_239_dout[15]),
  .I1(rom16_inst_255_dout[15]),
  .S0(ad[4])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_225),
  .I1(mux_o_226),
  .S0(ad[5])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_227),
  .I1(mux_o_228),
  .S0(ad[5])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_229),
  .I1(mux_o_230),
  .S0(ad[5])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_231),
  .I1(mux_o_232),
  .S0(ad[5])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(ad[6])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(ad[6])
);
MUX2 mux_inst_239 (
  .O(dout[15]),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(ad[7])
);
endmodule //Gowin_ROM16
