//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Thu Apr 07 21:09:13 2022

module Gowin_rPLL (clkout, clkoutd, clkin);

    output clkout;
    output clkoutd;
    input clkin;

    wire lock_o;
    wire clkoutp_o;
    wire clkoutd3_o;
    wire gw_gnd;

    assign gw_gnd = 1'b0;

    rPLL rpll_inst (
             .CLKOUT(clkout),
             .LOCK(lock_o),
             .CLKOUTP(clkoutp_o),
             .CLKOUTD(clkoutd),
             .CLKOUTD3(clkoutd3_o),
             .RESET(gw_gnd),
             .RESET_P(gw_gnd),
             .CLKIN(clkin),
             .CLKFB(gw_gnd),
             .FBDSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
             .IDSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
             .ODSEL({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
             .PSDA({gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
             .DUTYDA({gw_gnd,gw_gnd,gw_gnd,gw_gnd}),
             .FDLY({gw_gnd,gw_gnd,gw_gnd,gw_gnd})
         );

    defparam rpll_inst.FCLKIN = "27";
    defparam rpll_inst.DYN_IDIV_SEL = "false";
    defparam rpll_inst.IDIV_SEL = 2;
    defparam rpll_inst.DYN_FBDIV_SEL = "false";
    defparam rpll_inst.FBDIV_SEL = 7;
    defparam rpll_inst.DYN_ODIV_SEL = "false";
    defparam rpll_inst.ODIV_SEL = 8;
    defparam rpll_inst.PSDA_SEL = "0000";
    defparam rpll_inst.DYN_DA_EN = "true";
    defparam rpll_inst.DUTYDA_SEL = "1000";
    defparam rpll_inst.CLKOUT_FT_DIR = 1'b1;
    defparam rpll_inst.CLKOUTP_FT_DIR = 1'b1;
    defparam rpll_inst.CLKOUT_DLY_STEP = 0;
    defparam rpll_inst.CLKOUTP_DLY_STEP = 0;
    defparam rpll_inst.CLKFB_SEL = "internal";
    defparam rpll_inst.CLKOUT_BYPASS = "false";
    defparam rpll_inst.CLKOUTP_BYPASS = "false";
    defparam rpll_inst.CLKOUTD_BYPASS = "false";
    defparam rpll_inst.DYN_SDIV_SEL = 2;
    defparam rpll_inst.CLKOUTD_SRC = "CLKOUT";
    defparam rpll_inst.CLKOUTD3_SRC = "CLKOUT";
    defparam rpll_inst.DEVICE = "GW1NR-9C";

endmodule //Gowin_rPLL
