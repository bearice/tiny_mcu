//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NR-LV9QN88C6/I5
//Device: GW1NR-9C
//Created Time: Thu Apr 07 21:09:13 2022

module VRam (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [15:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [11:0] ada;
input [15:0] din;
input [11:0] adb;

wire [23:0] sdpb_inst_0_dout_w;
wire [7:0] sdpb_inst_0_dout;
wire [23:0] sdpb_inst_1_dout_w;
wire [15:8] sdpb_inst_1_dout;
wire [15:0] sdpb_inst_2_dout_w;
wire [15:0] sdpb_inst_2_dout;
wire dff_q_0;
wire gw_vcc;
wire gw_gnd;

assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[23:0],sdpb_inst_0_dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[11]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 8;
defparam sdpb_inst_0.BIT_WIDTH_1 = 8;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_0B = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_19 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_1A = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_1B = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_1C = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_1D = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_1E = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_1F = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_20 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_21 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_22 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_23 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_24 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_25 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_26 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_27 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_28 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_29 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_2A = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_2B = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_2C = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_2D = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_2E = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_2F = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_30 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_31 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_32 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_33 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_34 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_35 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_36 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_37 = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_38 = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_39 = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_3A = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_3B = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_3C = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;
defparam sdpb_inst_0.INIT_RAM_3D = 256'h6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C654821646C72;
defparam sdpb_inst_0.INIT_RAM_3E = 256'h21646C726F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F;
defparam sdpb_inst_0.INIT_RAM_3F = 256'h6F57206F6C6C654821646C726F57206F6C6C654821646C726F57206F6C6C6548;

SDPB sdpb_inst_1 (
    .DO({sdpb_inst_1_dout_w[23:0],sdpb_inst_1_dout[15:8]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,ada[11]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[11]}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:8]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_1.READ_MODE = 1'b0;
defparam sdpb_inst_1.BIT_WIDTH_0 = 8;
defparam sdpb_inst_1.BIT_WIDTH_1 = 8;
defparam sdpb_inst_1.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_1.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_1.RESET_MODE = "SYNC";
defparam sdpb_inst_1.INIT_RAM_00 = 256'h101F1E1D1C1B1A1908070605040302010F0E0D0CFBFAF9F8F7F6F5F4F3F2F1F0;
defparam sdpb_inst_1.INIT_RAM_01 = 256'h4241404F3E3D3C3B3A3938373635343221202F2E2D2C2B2A2928272615141312;
defparam sdpb_inst_1.INIT_RAM_02 = 256'h64636261606F6E6D6C6B6A6958575654535251505F5E5D5C4B4A494847464543;
defparam sdpb_inst_1.INIT_RAM_03 = 256'h969594939291909F8E8D8C8B8A8987868584838271707F7E7D7C7B7A79787675;
defparam sdpb_inst_1.INIT_RAM_04 = 256'hC8C7C6C5B4B3B2B1B0BFBEBDBCBAB9B8A7A6A5A4A3A2A1A0AFAEADAC9B9A9897;
defparam sdpb_inst_1.INIT_RAM_05 = 256'hEAE9E8E7E6E5E4E3E2E1E0EFDEDCDBDAD9D8D7D6D5D4D3D2C1C0CFCECDCBCAC9;
defparam sdpb_inst_1.INIT_RAM_06 = 256'h1C1B1A1918171615040302010F0E0D0C0B0A0908F7F6F5F4F3F2F1F0FEFDFCFB;
defparam sdpb_inst_1.INIT_RAM_07 = 256'h4E4D4C4B3A3938373635343231303F3E2D2C2B2A2928272625242321101F1E1D;
defparam sdpb_inst_1.INIT_RAM_08 = 256'h606F6E6D6C6B6A6968676564535251505F5E5D5C5B5A5958474645434241404F;
defparam sdpb_inst_1.INIT_RAM_09 = 256'h9291909F9E9D9C9B8A8987868584838281808F8E7D7C7B7A7978767574737271;
defparam sdpb_inst_1.INIT_RAM_0A = 256'hC4C3C2C1B0BFBEBDBCBAB9B8B7B6B5B4A3A2A1A0AFAEADACABA9A8A796959493;
defparam sdpb_inst_1.INIT_RAM_0B = 256'hE6E5E4E3E2E1E0EFEDECEBEAD9D8D7D6D5D4D3D2D1D0DFDECDCBCAC9C8C7C6C5;
defparam sdpb_inst_1.INIT_RAM_0C = 256'h18171615141312100F0E0D0C0B0A090807060504F3F2F1F0FEFDFCFBFAF9F8F7;
defparam sdpb_inst_1.INIT_RAM_0D = 256'h4A4948473635343231303F3E3D3C3B3A2928272625242321202F2E2D1C1B1A19;
defparam sdpb_inst_1.INIT_RAM_0E = 256'h6C6B6A6968676564636261605F5E5D5C5B5A5958575654534241404F4E4D4C4B;
defparam sdpb_inst_1.INIT_RAM_0F = 256'h9E9D9C9B9A9897968584838281808F8E8D8C8B8A7978767574737271707F7E7D;
defparam sdpb_inst_1.INIT_RAM_10 = 256'hC0CFCECDBCBAB9B8B7B6B5B4B3B2B1B0AFAEADACABA9A8A7A6A5A4A39291909F;
defparam sdpb_inst_1.INIT_RAM_11 = 256'hE2E1E0EFEDECEBEAE9E8E7E6D5D4D3D2D1D0DFDEDCDBDAD9C8C7C6C5C4C3C2C1;
defparam sdpb_inst_1.INIT_RAM_12 = 256'h141312101F1E1D1C0B0A0908070605040302010FFEFDFCFBFAF9F8F7F6F5F4F3;
defparam sdpb_inst_1.INIT_RAM_13 = 256'h4645434231303F3E3D3C3B3A3938373625242321202F2E2D2C2B2A2918171615;
defparam sdpb_inst_1.INIT_RAM_14 = 256'h68676564636261606F6E6D6C5B5A5958575654535251505F4E4D4C4B4A494847;
defparam sdpb_inst_1.INIT_RAM_15 = 256'h9A9897969594939281808F8E8D8C8B8A8987868574737271707F7E7D7C7B7A79;
defparam sdpb_inst_1.INIT_RAM_16 = 256'hCBCAC9C8B7B6B5B4B3B2B1B0BFBEBDBCABA9A8A7A6A5A4A3A2A1A0AF9E9D9C9B;
defparam sdpb_inst_1.INIT_RAM_17 = 256'hEDECEBEAE9E8E7E6E5E4E3E2D1D0DFDEDCDBDAD9D8D7D6D5C4C3C2C1C0CFCECD;
defparam sdpb_inst_1.INIT_RAM_18 = 256'h1F1E1D1C1B1A1918070605040302010F0E0D0C0BFAF9F8F7F6F5F4F3F2F1F0FE;
defparam sdpb_inst_1.INIT_RAM_19 = 256'h41404F4E3D3C3B3A3938373635343231202F2E2D2C2B2A292827262514131210;
defparam sdpb_inst_1.INIT_RAM_1A = 256'h636261606F6E6D6C6B6A6968575654535251505F5E5D5C5B4A49484746454342;
defparam sdpb_inst_1.INIT_RAM_1B = 256'h9594939291909F9E8D8C8B8A8987868584838281707F7E7D7C7B7A7978767574;
defparam sdpb_inst_1.INIT_RAM_1C = 256'hC7C6C5C4B3B2B1B0BFBEBDBCBAB9B8B7A6A5A4A3A2A1A0AFAEADACAB9A989796;
defparam sdpb_inst_1.INIT_RAM_1D = 256'hE9E8E7E6E5E4E3E2E1E0EFEDDCDBDAD9D8D7D6D5D4D3D2D1C0CFCECDCBCAC9C8;
defparam sdpb_inst_1.INIT_RAM_1E = 256'h1B1A1918171615140302010F0E0D0C0B0A090807F6F5F4F3F2F1F0FEFDFCFBFA;
defparam sdpb_inst_1.INIT_RAM_1F = 256'h4D4C4B4A3938373635343231303F3E3D2C2B2A2928272625242321201F1E1D1C;
defparam sdpb_inst_1.INIT_RAM_20 = 256'h6F6E6D6C6B6A6968676564635251505F5E5D5C5B5A5958574645434241404F4E;
defparam sdpb_inst_1.INIT_RAM_21 = 256'h91909F9E9D9C9B9A8987868584838281808F8E8D7C7B7A797876757473727170;
defparam sdpb_inst_1.INIT_RAM_22 = 256'hC3C2C1C0BFBEBDBCBAB9B8B7B6B5B4B3A2A1A0AFAEADACABA9A8A7A695949392;
defparam sdpb_inst_1.INIT_RAM_23 = 256'hE5E4E3E2E1E0EFEDECEBEAE9D8D7D6D5D4D3D2D1D0DFDEDCCBCAC9C8C7C6C5C4;
defparam sdpb_inst_1.INIT_RAM_24 = 256'h171615141312101F0E0D0C0B0A09080706050403F2F1F0FEFDFCFBFAF9F8F7F6;
defparam sdpb_inst_1.INIT_RAM_25 = 256'h4948474635343231303F3E3D3C3B3A3928272625242321202F2E2D2C1B1A1918;
defparam sdpb_inst_1.INIT_RAM_26 = 256'h6B6A6968676564636261606F5E5D5C5B5A5958575654535241404F4E4D4C4B4A;
defparam sdpb_inst_1.INIT_RAM_27 = 256'h9D9C9B9A9897969584838281808F8E8D8C8B8A8978767574737271707F7E7D7C;
defparam sdpb_inst_1.INIT_RAM_28 = 256'hCFCECDCBBAB9B8B7B6B5B4B3B2B1B0BFAEADACABA9A8A7A6A5A4A3A291909F9E;
defparam sdpb_inst_1.INIT_RAM_29 = 256'hE1E0EFEDECEBEAE9E8E7E6E5D4D3D2D1D0DFDEDCDBDAD9D8C7C6C5C4C3C2C1C0;
defparam sdpb_inst_1.INIT_RAM_2A = 256'h1312101F1E1D1C1B0A0908070605040302010F0EFDFCFBFAF9F8F7F6F5F4F3F2;
defparam sdpb_inst_1.INIT_RAM_2B = 256'h45434241303F3E3D3C3B3A3938373635242321202F2E2D2C2B2A292817161514;
defparam sdpb_inst_1.INIT_RAM_2C = 256'h676564636261606F6E6D6C6B5A5958575654535251505F5E4D4C4B4A49484746;
defparam sdpb_inst_1.INIT_RAM_2D = 256'h9897969594939291808F8E8D8C8B8A8987868584737271707F7E7D7C7B7A7978;
defparam sdpb_inst_1.INIT_RAM_2E = 256'hCAC9C8C7B6B5B4B3B2B1B0BFBEBDBCBAA9A8A7A6A5A4A3A2A1A0AFAE9D9C9B9A;
defparam sdpb_inst_1.INIT_RAM_2F = 256'hECEBEAE9E8E7E6E5E4E3E2E1D0DFDEDCDBDAD9D8D7D6D5D4C3C2C1C0CFCECDCB;
defparam sdpb_inst_1.INIT_RAM_30 = 256'h1E1D1C1B1A1918170605040302010F0E0D0C0B0AF9F8F7F6F5F4F3F2F1F0FEFD;
defparam sdpb_inst_1.INIT_RAM_31 = 256'h404F4E4D3C3B3A3938373635343231302F2E2D2C2B2A2928272625241312101F;
defparam sdpb_inst_1.INIT_RAM_32 = 256'h6261606F6E6D6C6B6A6968675654535251505F5E5D5C5B5A4948474645434241;
defparam sdpb_inst_1.INIT_RAM_33 = 256'h94939291909F9E9D8C8B8A8987868584838281807F7E7D7C7B7A797876757473;
defparam sdpb_inst_1.INIT_RAM_34 = 256'hC6C5C4C3B2B1B0BFBEBDBCBAB9B8B7B6A5A4A3A2A1A0AFAEADACABA998979695;
defparam sdpb_inst_1.INIT_RAM_35 = 256'hE8E7E6E5E4E3E2E1E0EFEDECDBDAD9D8D7D6D5D4D3D2D1D0CFCECDCBCAC9C8C7;
defparam sdpb_inst_1.INIT_RAM_36 = 256'h1A1918171615141302010F0E0D0C0B0A09080706F5F4F3F2F1F0FEFDFCFBFAF9;
defparam sdpb_inst_1.INIT_RAM_37 = 256'h4C4B4A4938373635343231303F3E3D3C2B2A2928272625242321202F1E1D1C1B;
defparam sdpb_inst_1.INIT_RAM_38 = 256'h6E6D6C6B6A6968676564636251505F5E5D5C5B5A5958575645434241404F4E4D;
defparam sdpb_inst_1.INIT_RAM_39 = 256'h909F9E9D9C9B9A9887868584838281808F8E8D8C7B7A7978767574737271707F;
defparam sdpb_inst_1.INIT_RAM_3A = 256'hC2C1C0CFBEBDBCBAB9B8B7B6B5B4B3B2A1A0AFAEADACABA9A8A7A6A594939291;
defparam sdpb_inst_1.INIT_RAM_3B = 256'hE4E3E2E1E0EFEDECEBEAE9E8D7D6D5D4D3D2D1D0DFDEDCDBCAC9C8C7C6C5C4C3;
defparam sdpb_inst_1.INIT_RAM_3C = 256'h1615141312101F1E0D0C0B0A0908070605040302F1F0FEFDFCFBFAF9F8F7F6F5;
defparam sdpb_inst_1.INIT_RAM_3D = 256'h48474645343231303F3E3D3C3B3A3938272625242321202F2E2D2C2B1A191817;
defparam sdpb_inst_1.INIT_RAM_3E = 256'h6A6968676564636261606F6E5D5C5B5A5958575654535251404F4E4D4C4B4A49;
defparam sdpb_inst_1.INIT_RAM_3F = 256'h9C9B9A9897969594838281808F8E8D8C8B8A8987767574737271707F7E7D7C7B;

SDPB sdpb_inst_2 (
    .DO({sdpb_inst_2_dout_w[15:0],sdpb_inst_2_dout[15:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,ada[11],ada[10]}),
    .BLKSELB({gw_gnd,adb[11],adb[10]}),
    .ADA({ada[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]}),
    .ADB({adb[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_2.READ_MODE = 1'b0;
defparam sdpb_inst_2.BIT_WIDTH_0 = 16;
defparam sdpb_inst_2.BIT_WIDTH_1 = 16;
defparam sdpb_inst_2.BLK_SEL_0 = 3'b010;
defparam sdpb_inst_2.BLK_SEL_1 = 3'b010;
defparam sdpb_inst_2.RESET_MODE = "SYNC";
defparam sdpb_inst_2.INIT_RAM_00 = 256'hAD21AC64AB6CA972A86FA757A620A56FA46CA36CA265A14890219F649E6C9D72;
defparam sdpb_inst_2.INIT_RAM_01 = 256'hCE6CCD6CCB65CA48B921B864B76CB672B56FB457B320B26FB16CB06CBF65BE48;
defparam sdpb_inst_2.INIT_RAM_02 = 256'hDF6FDE57DC20DB6FDA6CD96CD865D748C621C564C46CC372C26FC157C020CF6F;
defparam sdpb_inst_2.INIT_RAM_03 = 256'hE021EF64ED6CEC72EB6FEA57E920E86FE76CE66CE565E448D321D264D16CD072;
defparam sdpb_inst_2.INIT_RAM_04 = 256'h016C0F6C0E650D48FC21FB64FA6CF972F86FF757F620F56FF46CF36CF265F148;
defparam sdpb_inst_2.INIT_RAM_05 = 256'h126F10571F201E6F1D6C1C6C1B651A4809210864076C0672056F04570320026F;
defparam sdpb_inst_2.INIT_RAM_06 = 256'h23212164206C2F722E6F2D572C202B6F2A6C296C2865274816211564146C1372;
defparam sdpb_inst_2.INIT_RAM_07 = 256'h436C426C416540483F213E643D6C3C723B6F3A573920386F376C366C35653448;
defparam sdpb_inst_2.INIT_RAM_08 = 256'h546F53575220516F506C5F6C5E655D484C214B644A6C4972486F47574620456F;
defparam sdpb_inst_2.INIT_RAM_09 = 256'h65216464636C6272616F60576F206E6F6D6C6C6C6B656A4859215864576C5672;
defparam sdpb_inst_2.INIT_RAM_0A = 256'h866C856C8465834872217164706C7F727E6F7D577C207B6F7A6C796C78657648;
defparam sdpb_inst_2.INIT_RAM_0B = 256'h976F96579520946F936C926C916590488F218E648D6C8C728B6F8A578920876F;
defparam sdpb_inst_2.INIT_RAM_0C = 256'hA821A764A66CA572A46FA357A220A16FA06CAF6CAE65AD489C219B649A6C9872;
defparam sdpb_inst_2.INIT_RAM_0D = 256'hC96CC86CC765C648B521B464B36CB272B16FB057BF20BE6FBD6CBC6CBA65B948;
defparam sdpb_inst_2.INIT_RAM_0E = 256'hDA6FD957D820D76FD66CD56CD465D348C221C164C06CCF72CE6FCD57CB20CA6F;
defparam sdpb_inst_2.INIT_RAM_0F = 256'hEB21EA64E96CE872E76FE657E520E46FE36CE26CE165E048DF21DE64DC6CDB72;
defparam sdpb_inst_2.INIT_RAM_10 = 256'h0C6C0B6C0A650948F821F764F66CF572F46FF357F220F16FF06CFE6CFD65FC48;
defparam sdpb_inst_2.INIT_RAM_11 = 256'h1D6F1C571B201A6F196C186C1765164805210464036C0272016F0F570E200D6F;
defparam sdpb_inst_2.INIT_RAM_12 = 256'h2E212D642C6C2B722A6F29572820276F266C256C24652348122110641F6C1E72;
defparam sdpb_inst_2.INIT_RAM_13 = 256'h4F6C4E6C4D654C483B213A64396C3872376F36573520346F326C316C30653F48;
defparam sdpb_inst_2.INIT_RAM_14 = 256'h506F5F575E205D6F5C6C5B6C5A65594848214764466C4572436F42574120406F;
defparam sdpb_inst_2.INIT_RAM_15 = 256'h612160646F6C6E726D6F6C576B206A6F696C686C6765654854215364526C5172;
defparam sdpb_inst_2.INIT_RAM_16 = 256'h826C816C80658F487E217D647C6C7B727A6F79577820766F756C746C73657248;
defparam sdpb_inst_2.INIT_RAM_17 = 256'h936F92579120906F9F6C9E6C9D659C488B218A64896C8772866F85578420836F;
defparam sdpb_inst_2.INIT_RAM_18 = 256'hA421A364A26CA172A06FAF57AE20AD6FAC6CAB6CA965A84897219664956C9472;
defparam sdpb_inst_2.INIT_RAM_19 = 256'hC56CC46CC365C248B121B064BF6CBE72BD6FBC57BA20B96FB86CB76CB665B548;
defparam sdpb_inst_2.INIT_RAM_1A = 256'hD66FD557D420D36FD26CD16CD065DF48CE21CD64CB6CCA72C96FC857C720C66F;
defparam sdpb_inst_2.INIT_RAM_1B = 256'hE721E664E56CE472E36FE257E120E06FEF6CED6CEC65EB48DA21D964D86CD772;
defparam sdpb_inst_2.INIT_RAM_1C = 256'h086C076C06650548F421F364F26CF172F06FFE57FD20FC6FFB6CFA6CF965F848;
defparam sdpb_inst_2.INIT_RAM_1D = 256'h196F18571720166F156C146C1365124801210F640E6C0D720C6F0B570A20096F;
defparam sdpb_inst_2.INIT_RAM_1E = 256'h2A212964286C2772266F25572420236F216C206C2F652E481D211C641B6C1A72;
defparam sdpb_inst_2.INIT_RAM_1F = 256'h4B6C4A6C4965484837213664356C3472326F315730203F6F3E6C3D6C3C653B48;
defparam sdpb_inst_2.INIT_RAM_20 = 256'h5C6F5B575A20596F586C576C5665544843214264416C40724F6F4E574D204C6F;
defparam sdpb_inst_2.INIT_RAM_21 = 256'h6D216C646B6C6A72696F68576720656F646C636C6265614850215F645E6C5D72;
defparam sdpb_inst_2.INIT_RAM_22 = 256'h8E6C8D6C8C658B487A217964786C7672756F74577320726F716C706C7F657E48;
defparam sdpb_inst_2.INIT_RAM_23 = 256'h9F6F9E579D209C6F9B6C9A6C9865974886218564846C8372826F815780208F6F;
defparam sdpb_inst_2.INIT_RAM_24 = 256'hA021AF64AE6CAD72AC6FAB57A920A86FA76CA66CA565A44893219264916C9072;
defparam sdpb_inst_2.INIT_RAM_25 = 256'hC16CC06CCF65CE48BD21BC64BA6CB972B86FB757B620B56FB46CB36CB265B148;
defparam sdpb_inst_2.INIT_RAM_26 = 256'hD26FD157D020DF6FDE6CDC6CDB65DA48C921C864C76CC672C56FC457C320C26F;
defparam sdpb_inst_2.INIT_RAM_27 = 256'hE321E264E16CE072EF6FED57EC20EB6FEA6CE96CE865E748D621D564D46CD372;
defparam sdpb_inst_2.INIT_RAM_28 = 256'h046C036C02650148F021FE64FD6CFC72FB6FFA57F920F86FF76CF66CF565F448;
defparam sdpb_inst_2.INIT_RAM_29 = 256'h156F14571320126F106C1F6C1E651D480C210B640A6C0972086F07570620056F;
defparam sdpb_inst_2.INIT_RAM_2A = 256'h26212564246C2372216F20572F202E6F2D6C2C6C2B652A4819211864176C1672;
defparam sdpb_inst_2.INIT_RAM_2B = 256'h476C466C4565434832213164306C3F723E6F3D573C203B6F3A6C396C38653748;
defparam sdpb_inst_2.INIT_RAM_2C = 256'h586F57575620546F536C526C516550484F214E644D6C4C724B6F4A574920486F;
defparam sdpb_inst_2.INIT_RAM_2D = 256'h69216864676C6572646F63576220616F606C6F6C6E656D485C215B645A6C5972;
defparam sdpb_inst_2.INIT_RAM_2E = 256'h8A6C896C8765864875217464736C7272716F70577F207E6F7D6C7C6C7B657A48;
defparam sdpb_inst_2.INIT_RAM_2F = 256'h9B6F9A579820976F966C956C9465934882218164806C8F728E6F8D578C208B6F;
defparam sdpb_inst_2.INIT_RAM_30 = 256'hAC21AB64A96CA872A76FA657A520A46FA36CA26CA165A0489F219E649D6C9C72;
defparam sdpb_inst_2.INIT_RAM_31 = 256'hCD6CCB6CCA65C948B821B764B66CB572B46FB357B220B16FB06CBF6CBE65BD48;
defparam sdpb_inst_2.INIT_RAM_32 = 256'hDE6FDC57DB20DA6FD96CD86CD765D648C521C464C36CC272C16FC057CF20CE6F;
defparam sdpb_inst_2.INIT_RAM_33 = 256'hEF21ED64EC6CEB72EA6FE957E820E76FE66CE56CE465E348D221D164D06CDF72;
defparam sdpb_inst_2.INIT_RAM_34 = 256'h0F6C0E6C0D650C48FB21FA64F96CF872F76FF657F520F46FF36CF26CF165F048;
defparam sdpb_inst_2.INIT_RAM_35 = 256'h106F1F571E201D6F1C6C1B6C1A65194808210764066C0572046F03570220016F;
defparam sdpb_inst_2.INIT_RAM_36 = 256'h212120642F6C2E722D6F2C572B202A6F296C286C2765264815211464136C1272;
defparam sdpb_inst_2.INIT_RAM_37 = 256'h426C416C40654F483E213D643C6C3B723A6F39573820376F366C356C34653248;
defparam sdpb_inst_2.INIT_RAM_38 = 256'h536F52575120506F5F6C5E6C5D655C484B214A64496C4872476F46574520436F;
defparam sdpb_inst_2.INIT_RAM_39 = 256'h64216364626C6172606F6F576E206D6F6C6C6B6C6A65694858215764566C5472;
defparam sdpb_inst_2.INIT_RAM_3A = 256'h856C846C83658248712170647F6C7E727D6F7C577B207A6F796C786C76657548;
defparam sdpb_inst_2.INIT_RAM_3B = 256'h000000000000000000000000000000008E218D648C6C8B728A6F89578720866F;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(adb[11]),
  .CLK(clkb),
  .CE(ceb)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(sdpb_inst_0_dout[0]),
  .I1(sdpb_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(sdpb_inst_0_dout[1]),
  .I1(sdpb_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(sdpb_inst_0_dout[2]),
  .I1(sdpb_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(sdpb_inst_0_dout[3]),
  .I1(sdpb_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(sdpb_inst_0_dout[4]),
  .I1(sdpb_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(sdpb_inst_0_dout[5]),
  .I1(sdpb_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(sdpb_inst_0_dout[6]),
  .I1(sdpb_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(sdpb_inst_0_dout[7]),
  .I1(sdpb_inst_2_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(dout[8]),
  .I0(sdpb_inst_1_dout[8]),
  .I1(sdpb_inst_2_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[9]),
  .I0(sdpb_inst_1_dout[9]),
  .I1(sdpb_inst_2_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(dout[10]),
  .I0(sdpb_inst_1_dout[10]),
  .I1(sdpb_inst_2_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(dout[11]),
  .I0(sdpb_inst_1_dout[11]),
  .I1(sdpb_inst_2_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_38 (
  .O(dout[12]),
  .I0(sdpb_inst_1_dout[12]),
  .I1(sdpb_inst_2_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_41 (
  .O(dout[13]),
  .I0(sdpb_inst_1_dout[13]),
  .I1(sdpb_inst_2_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(dout[14]),
  .I0(sdpb_inst_1_dout[14]),
  .I1(sdpb_inst_2_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_47 (
  .O(dout[15]),
  .I0(sdpb_inst_1_dout[15]),
  .I1(sdpb_inst_2_dout[15]),
  .S0(dff_q_0)
);
endmodule //VRam
