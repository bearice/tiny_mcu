//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NZ-LV1QN48C6/I5
//Device: GW1NZ-1
//Created Time: Sun Apr 03 21:48:52 2022

module FontRom (dout, clk, oce, ce, reset, ad);

output [0:0] dout;
input clk;
input oce;
input ce;
input reset;
input [13:0] ad;

wire [30:0] prom_inst_0_dout_w;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h000000384482BAC68282AA824438000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000010387CFEFEFEEE4400000000000000387CFEC6BAFEFED6FE7C380000;
defparam prom_inst_0.INIT_RAM_02 = 256'h000000007C10EEFED6383838000000000000000010387CFEFE7C381000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000000000183C3C18000000000000000000007C10D6FEFE7C381000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h00000000001824424224180000000000FFFFFFFFFFFFE7C3C3E7FFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000003C6666666666BCE0C0F080000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000C1C1C18101010D070301000000000000018187E18183C6666663C0000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000010927C44C6447C9210000000000060E6EECE8C88888888E8F8180000;
defparam prom_inst_0.INIT_RAM_08 = 256'h000000000030383C3E3C38300000000000000000000C1C3C7C3C1C0C00000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h000000666600666666666666666600000000000010387C101010107C38100000;
defparam prom_inst_0.INIT_RAM_0A = 256'h00007CC660386CC6C66C380CC67C00000000000090909090909C9E9E9EFC0000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000007C10387C101010107C3810000000000000000000FEFEFEFE0000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000010387C10101010101010000000000000101010101010107C38100000;
defparam prom_inst_0.INIT_RAM_0D = 256'h00000000000000080CFE0C0800000000000000000000002060FE602000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h000000000000002466FF662400000000000000000000FE060606060000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h00000000000010387CFEFE0000000000000000000000FEFE7C38100000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000001818001818181818181818000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h000000006C6CFE6C6C6CFE6C6C00000000000000000000000000666666660000;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000060F2660C183060CC9E0C00000010107CD6D0C07C0616D67C10100000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000000000000000000000181818180000000000DC666666D61C386C6C380000;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000C181830303030303018180C000000006030301818181818183030600000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000000018187E181800000000000000000000105438FE38541000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000000000007E0000000000000000000810181800000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000006060C0C181830306060000000000000181800000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000030303030303030303C300000000000007CC6C6C6C6D6C6C6C67C000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000003C66626060386060663C0000000000007E06060C18306066663C000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000003C66626060663E06067E0000000000006060FE6266646C687870000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000001818181830303060607E0000000000003C666666663E06060C38000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000001C3060607C666666663C0000000000003C666666663C2466663C000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000081018180000001818000000000000000000181800000018180000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000007C00007C000000000000000000006030180C060C183060000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h000018180018183060C0C6C67C000000000000000C183060C06030180C000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h000000C6C6C6C6FEC6C6C66C38000000000078CC06F6D6D6B6F6C6CC78000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000007CC6C606060606C6C67C0000000000007EC6C6C6C67EC6C6C67E000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h000000FE060606067E060606FE0000000000003E66C6C6C6C6C6C6663E000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h000000DCE6C6C6E60606C6C67C00000000000006060606067E060606FE000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000003C18181818181818183C000000000000C6C6C6C6C6FEC6C6C6C6000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h000000C6C666361E1E3666C6C60000000000003C6666606060606060F8000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h000000C6C6C6C6D6D6FEEEC682000000000000FE060606060606060606000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000007CC6C6C6C6C6C6C6C67C000000000000C6C6C6C6E6F6DECEC6C2000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h00E0307CC6C6C6C6C6C6C6C67C000000000000060606067EC6C6C6C67E000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000007CC6C6E0701C0EC6C67C000000000000C6C666367EC6C6C6C67E000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000007CC6C6C6C6C6C6C6C6C60000000000001818181818181818187E000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000006C6CD6D6D6C6C6C6C6C600000000000038386C6CC6C6C6C6C6C6000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h00000018181818183C66666666000000000000C6C6C66C38386CC6C6C6000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h00007818181818181818181818780000000000FE0C0C181830306060FE000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h00003C303030303030303030303C00000000006060303018180C0C0606000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h00FF000000000000000000000000000000000000000000000000C66C38100000;
defparam prom_inst_0.INIT_RAM_30 = 256'h000000FCC6C6FCC0C07C000000000000000000000000000000000030180C0000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000007CC6060606C67C0000000000000000007EC6C6C6C6CE76060606000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000007C0606FEC6C67C000000000000000000FCC6C6C6C6E6DCC0C0C0000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h007CC0C0DCE6C6C6C6FC0000000000000000001818181818187E1818F0000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h000000FC30303030303C003030000000000000C6C6C6C6C6CE76060606000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h000000C666361E1E3666060606000000001E30303030303030303C0030300000;
defparam prom_inst_0.INIT_RAM_36 = 256'h000000C6C6D6D6D6FE6E0000000000000000007018181818181818181C000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000007CC6C6C6C6C67C000000000000000000C6C6C6C6C6CE76000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h00C0C0C0DCE6C6C6C6FC000000000000000606067EC6C6C6CE76000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000007CC6C07C06C67C0000000000000000000C0C0C0C0CDC6C000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h000000DCE6C6C6C6C6C60000000000000000007018181818187E181810000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000006C7CD6D6D6C6C600000000000000000038386C6CC6C6C6000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h007CC0C0DCE6C6C6C6C6000000000000000000C6C66C386CC6C6000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h007018181818180E1818181818700000000000FE060C183060FE000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h001C3030303030E030303030301C000000181818181818181818181818181800;
defparam prom_inst_0.INIT_RAM_3F = 256'h00000000FE828282C66C381000000000000000000000000000000062FE8C0000;

endmodule //FontRom
